Vad fan ? Typiskt . 
Hej . 
Jag ... Jag såg din jobbannons . 
LAGERARBETE OCH ENKLA UPPGIFTER Jag är Jeongmin Bae . 
Vi har träffats . 
Jag gick i skolan med Jian . 
Hur funkar den ? 
Jag pratade inte med dig . 
Hur många gånger måste jag säga det ? 
Jag var nära att dö . 
Hur som helst , jag är inne . 
Du såg väl bilden på Jian ? 
Du får murthehelps källa senare idag . 
Du fick varuhuset på tre dagar . Det är tack vare mig . 
Va ? 
Ska jag döda henne ? 
Vadå ? 
Kan du inte avsluta jobbet ? 
Kan du inte bättre ? 
Vad menade du ? Låste du in mig ? 
Va ? 
Det du sa innan . 
Att när vi var små så låste du in mig i skolförrådet . 
Jaha , det ... 
Jinman Jeong ! 
Jinman Jeong ! 
För att se om du var stum på riktigt . 
Jag bad mina vänner göra det . 
Jag trodde att du kunde tala i kris . 
Du borde tacka mig . 
Du övervann din afasi . 
Du är nog förvirrad . 
Du vet inte vad som pågår . 
Det här var omöjligt att förutse , så jag förstår . 
Vad fan snackar du om ? 
Vill du veta ? Vad som händer just nu . 
Babylon existerar . 
Din idiot . 
Det finns inga lönnmördare här . 
Du såg ju sajten på mörka webben . 
Det var en vapenhandel . 
En AK-47 för 1,2 miljoner won . 
Vill du köpa en eller ? 
Du blev utkastad från militären , vad ska du med den till ? 
Kan du ens hantera en pistol ? 
Jösses . Har du någon koll alls ? 
Den här sajten var annorlunda . 
De återställde den på fem minuter . 
Det är ganska skumt . 
Lägg av ! 
Hög kvalitet betyder att det är fejk . 
Är du en amatör , eller ? 
Jag , amatör ? 
Vem är proffs då ? 
Vår högskola är okänd . Vi är inga proffs . 
Vi är nollor . 
Så många hackare försöker få drömjobb på stora företag . 
Alla äkta black hats i landet har gett upp . 
De har alla blivit white hat . 
Jag ska visa vad en black hat hackare är . 
Du kommer att hamna i fängelse . 
Är du rädd för fängelse ? 
Självklart ! 
- Så rädd ! - Sluta . 
Håll dig till dina grillspett . 
Vad är fel med det ? 
ANGE KOD Vad hette sidan ? 
Murthehelp . 
Jäklar . 
Vem fan röker inomhus nuförtiden ? 
Idioten blängde på oss . 
Ska vi spöa honom ? 
Han behöver nog en omgång . 
Jag har inte känt mig ... 
Hackade ni murthehelp ? 
En minut kvar . 
Det här är vansinne . 
Jag gjorde det ! 
Vänta . Jag klarar det ! Ge mig bara lite mer tid ! Jag är nästan klar ... 
En fråga ... Tar ni hand om kroppen ? 
Det var då jag insåg att jag var annorlunda . 
Berätta om min farbror , inte dig själv . 
Men allt hänger ihop . 
Ha lite tålamod . 
Känner du honom ? 
Hon då ? 
Förlåt . 
Jag var inte så här i militären . 
Jag har inte tränat sen jag kom hem . 
Vila en stund . 
Okej . 
Jag måste verkligen träna . 
Den är felvänd . 
Skit också . 
Vad är det här ? 
Fan vad varmt det är . 
Helvete . 
Jag måste duscha . Fan . 
Vad fan letar jag efter ? 
Va ? 
Det var inget . 
Något att dricka . 
Tack . 
Hur mår Jian ? 
Vi var nära vänner i lågstadiet . 
DU HAR EN DAG KVAR Fan också ... 
Chefen ? Jag måste på toa . 
Får jag använda toaletten i huset ? 
Tack . 
Vad letar du efter ? 
Hej . Skrämde jag dig ? 
För att slippa gå fram och tillbaka när Jian är hemma , installerade jag en högtalare . 
Jag kikade bara runt lite . 
- Förlåt . - Det är lugnt . 
Förresten , visst pluggar du IT ? 
Ja , IT . 
Vad bra . 
Jag tror att min dator är sönder . 
Kan du laga den åt mig ? 
Jag lägger på extra på lönen . 
Visst . 
SKANNING PÅGÅR ... Du har nog fått ett virus . 
Jag sparar alla filer och formaterar datorn . 
Okej , tack . 
Hur mycket vill du ha för besväret ? 
Ingenting . 
Jian och jag var nära vänner . 
- Så det ... - I vilken årskurs ? 
Förlåt ? 
Jag har aldrig träffat Jians vänner . 
När blev ni vänner ? 
Jo ... När vi var jättesmå . 
I tvåan . 
Hon var oförskämd och hade inga vänner . 
Jian kunde inte prata så bra på den tiden . 
Jag brukade hjälpa henne . 
Och jag vet inte om du minns , men hon blev inlåst i skolan ... 
Ja , just det . 
Jag bjuder på middag sen . 
Jag går och städar . Kom när du är klar . Okej . 
Det gör jag . 
Det var lätt . 
Fy fan , jag luktar gödsel . 
Vem hade kunnat tro det här ? 
När är det klart ? 
ÄR DU KLAR ? Jinman Jeong måste logga in först . 
Vilka idioter . 
Han är inne . 
Så där ja . 
Det fungerade . 
Vad är det här ? 
Helvete . 
Lyssna noga . 
Om du dödar mig så var allt förgäves . 
Jag designade det så . 
Det är jag , Yonghan . 
Du har stake , grabben . 
För att vara säker . 
Dödar du mig så återställs murthehelp och du kommer inte in . 
Bara jag kan komma in . 
Döda honom . 
Vänta lite ! 
Vänta . 
Du såg mig jobba . 
Jag är bra på det här . 
Jag är bra på att hacka . 
Vad vill du ha ? 
Jinman Jeong ? 
Eller vapnen ? 
Jag har en riktigt grym plan . 
Jag lyssnar . 
Och allt gick enligt planen . 
Så pinsamt . Varför börjar det här ? 
Vad fan ? 
Så den stammande idioten bluffade . 
Jag trodde att man kunde se något . 
Det säger ingenting om vad som hände . 
Är du inte nyfiken , Jian ? 
Titta noga hur jag dödade din farbror . 
Hjälp , farbror ! 
Jag vet inte var jag är ! 
Fan , släpp mig ! 
Hjälp , farbror ! 
Jag vet inte var jag är ! 
Om du dödar mig , kommer Jian ... Hjälp , farbror ! 
- att dödas av Babylon . - Var är jag ? 
Sätt ner mig medan jag frågar snällt ! 
Nu ! 
Helvete ! Hjälp , farbror ! 
Jag vet inte var jag är ! 
Jag gör som du säger . 
Låt Jian gå som du lovade . 
Ja , självklart . 
Förtroende är viktigt i den här branschen . 
Lossa mig nu . 
Pasin . Behåll pengarna . 
Jinman Jeong ! 
Sätt ner mig ! 
Din jävel ! Hörru ! Helvete . 
Be Babylon att hålla sitt löfte . 
Nicka om du förstår . 
Helvete . 
Ett konstverk , eller hur ? 
Hur fick du min röst ? 
Jag har aldrig sagt det där . 
Det är en deepfake . 
Jag kan göra en på mindre än tio minuter . 
Och närbutikschefen hjälpte till med röstinspelningen . 
Kolla . 
Jian Jeong är dum i huvudet 
Jian Jeong är dum i huvudet 
Och din farbror var så ... 
Den store Jinman var dum nog att gå på det och begå självmord . 
Nej ! 
Jag var lite rädd eftersom de mäktiga Babylon var så försiktiga . 
Men jag oroade mig i onödan . 
Det var för enkelt . 
Men det betyder att jag är skicklig . 
En så svår sak var enkel för mig . 
Därför blev jag utvald . 
Vad är det ? 
Du är bara deras springpojke . 
Pratar du om mig ? 
Babylon ? 
De kommer att döda dig så fort du går ut härifrån . 
Nej , vänta . 
Om du dödar mig så dödar den där kvinnan dig först . 
Klarar du dig ? 
Du . Gör mig inte förbannad . 
Babylon bad mig nyss att döda dig . 
Men du , minns du inte 
vad du sa till mig ? 
" Alla med en kod måste skydda kod grön . " 
Min farbror är död , jag är den enda kod grön . 
Jag vet inte allt om Jinman ... Men av allt att döma är det nog fler som kommer att skydda mig . 
Vad snackar du om ? 
Använd hjärnan om du har en . 
Ingen från Babylon är här . De bryr sig inte om du dör . 
De där drönarna försökte döda oss . 
Du är utbytbar för dem . 
Den enda kod grön sitter framför dig . 
Det är mig du bör göra en deal med , 
inte dem . 
Vem är du att läxa upp mig ? 
Skulle jag förhandla med dig ? 
Jinman Jeong är död . 
Tror du att Murthehelp är ditt nu ? 
Du visste ingenting för några timmar sen . 
Du . Titta där . 
De kan ta sina drönare och idioter och skjuta vilt . Men jag tog mig hit och fångade dig . Jag ! 
Just det . 
Du gnydde och kröp runt i hallen för det här . 
Du kissade nästan på dig . 
Du kom så här långt för att Babylon tvingade dig , fegis ! 
Vad pratar du om ? 
Bara rädda idioter väsnas som hyenor ! 
Som du och skitstövlarna däruppe ! 
Säg ett ord till . 
Jävla subba . 
Jian ? 
Jian Jeong ! 
Du blev väl inte stum igen ? 
Använd allt omkring dig i krislägen . 
Använd alla medel för att överleva . 
Jag ska försöka . 
Vad fan ? 
Jag dödade nästan Jian innan . Och nu ska hon inte dö ? 
Tänk om jag redan hade dödat henne ? 
Är detta det bästa du kan göra ? 
Din lilla ... 
Behövs ansiktsigenkänning nu ? Skämtar du med mig ? 
Varför är du så sen , din skit ? 
Hej ! 
Var det därför ? 
Jag ville ge dig den här , men det var svårt . 
- Här finns bara berg . - Din lille skit . 
Hata mig inte . 
Din farbror var inget helgon . 
Jinman Jeong dödade många människor . 
Och Jian . Världen vi lever i ... Det handlar inte om att vara god eller ond , utan stark eller svag . 
Jinman var högst upp i näringskedjan och dog av fällan jag gillrade . 
Alltså är jag starkare än Jinman . 
Tror du att du kan fly ... 
Helvete ! Allvarligt ? 
Jian . 
Fan ! 
Jian Jeong ! 
Snälla ! 
Jian . 
Jian ! 
Jian , vänta . Du kan inte mäta dig med Jinman . 
Jian ... 
Tänk igenom det här . 
Ställ dig på min sida . 
När jättar kolliderar , faller de som din farbror . 
De svaga måste veta sin plats och välja klokt . 
Din dummer . 
Ja , visst . 
Hur kunde du lämna Jian ensam ? 
Hon måste lösa problemen på egen hand . 
Det är så hon lär sig att överleva . 
Som chefen ville . 
Oroa dig inte . 
Jian Jeong är inte svag . 
De attackerar snart igen . 
Är det här allt ? 
Bara 12 kulor ? 
Efter det som hände med Bale sa chefen att en attack kan ske när som helst . 
För att kunna försvara oss då , byggde han om . 
Så ... 
Vad gör du ? 
Det är så uppfriskande . 
Precis vad jag behövde ! 
Det var inte nödvändigt . 
Jag har varit sugen på sötsaker på sistone . 
Har du sparat ? 
Att vara anställd suger nuförtiden . Jag tänkte starta eget , som du . 
Det sägs att kontoret är ett slagfält , men utanför är ett helvete . 
Det kan jag intyga . 
Eftersom jag är ensam nu betalar jag varje kula ur egen ficka . 
Det är för jävligt . 
När man är med Babylon är inget olagligt . 
Det är sant . 
Stanna så länge du kan . 
Det har du rätt i . Jag tänkte mig inte för . 
Jäklar alltså . 
Förresten , det verkar som om Minhye dödade Kim . 
Den förbannade kärringen . 
Jävlar . 
Du har trimmat bilen . Går den bra ? 
Jag köpte den begagnad . 
Den kör som en dröm . Och den är robust . 
De är här . 
" Bubblans biltvätt . " 
Det ser så billigt ut . Varför biltvätt ? 
Sover du ? 
Vad liten den är . 
Värmer den upp eller ? 
De här betyder problem . 
Acceptera inte dem . 
De kommer att stjäla våra jobb i framtiden . 
Den är inte så bra som jag trodde . Är den inte lite töntig ? 
Attack påbörjas . 
De kan stjäla våra jobb redan nu . 
Vad gör ni ? 
Okej . Grupp 2 , hör ni mig ? 
Döda inte Jian Jeong . Fånga henne levande . 
Men det gör inget om ni bryter en arm eller ett ben . 
Okej . Akta er för Minhye . 
Håll er vid liv ! 
På ytan ser det ut som ett vanligt hus , men allt är byggt för försvar . 
Utnyttjar vi det kan ingen komma in . 
Kuma . Skynda dig . 
Vi klarar oss , om vi inte träffas av en missil . 
Hur ska du stoppa den ? 
In här , Minhye ! 
Vi kan ta oss in tack vare dig . 
Svara för fan . 
Gå in . 
Måste han svära ? 
Vad fan är det här för jalusi ? Vänta . 
Hur kom ni in ? 
Är vi instängda ? Oroa dig inte . 
Var inte rädda . 
Var inte rädda . 
När fixade Jinman det här ? 
Så klart att du inte kunde göra det lätt för oss . 
Din jävel . 
Gör något åt det där . 
Ska ni inte göra någonting ? 
De gömmer sig . 
Jinman tog inte hit mig för ett enkelt uppdrag . 
Du får klara dig själv nu . 
Vad vill du att jag ska göra ? 
Jian , du måste vara förvirrad . 
Vi har ont om tid men du måste välja . 
Ett . Om du vill fly från situationen gå till sidan 87 . 
Murthehelps bakdörr leder till en flyktväg . 
I slutet av den finns en ny identitet , pengar till ditt nya liv och telefonnumret till en person som kan hjälpa dig att börja om . 
Du får en ny identitet . 
Du kan glömma det här livet och börja om . 
Två . Om du vill kämpa med dina försvarare och de som kommer att stå vid din sida 
och att skydda denna plats , vänd bladet och läs guiden noggrant . 
Förlåt att du drogs in i detta kaos , men valet är ditt , Jian . 
Vad fan ... 
Det är gas ! Gas ! - Det är gas ! Gas ! - Gas ! 
Det här är självmord . 
Nu ! 
Var på er vakt . 
Minhye ! Här borta ! 
Helvete . 
Vad i helvete ? 
Vad var det ? 
En explosion ? 
Är du okej ? 
Har du fler kläder ? 
Minhye ! - Minhye ! - Så du är Jian Jeong . 
Släpp mig ! 
Släpp mig ! 
Och nu då ? 
Du är verkligen lik din farbror . 
Vad har du gjort med mitt ansikte ? 
Kuma , vad hände ? 
Har du Jian och Minhye ? 
Ja , jag har dem , men ... 
Alla andra är döda . 
Döda inte Jian än . 
Uppfattat . 
Jag skär bort halva ansiktet . 
Hon måste kännas igen . 
Mäster ? 
Vi har ont om tid . 
Gör dig redo . 
Bale är på väg . 
" Bale ? " 
Dina föräldrars mördare . 
Vad var det ? 
En slangbella ? 
Ni två får lösa det här . 
