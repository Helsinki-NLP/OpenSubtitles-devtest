Den nya inrikesministern är ung . 
Choi Minkyu . 
President Rhee favoriserar honom . 
Ska vi boka ett möte ? 
Minchul ordnar det . 
Hur var ritten ? 
Han är bra . Låt mig få honom . 
Ursäkta ? 
Du får min valkrets i utbyte mot den . 
Jag är fäst vid honom . 
Jag litar inte på nån politiker . 
Jag ska se till att du får en plats . 
Tack , allihop . 
Jag kom in i Nationalförsamlingen tack vare Cheongwooförbundet . 
Jag ska göra mitt bästa för er . 
När industrikomplexet är klart är Korea så gott som vårt . 
Vad sa Choi Minkyu ? 
Han ska prata med president Rhee och meddelar oss . 
Bad han om pengar ? 
Ja . 
Hur mycket pengar ska han roffa åt sig ? 
Be medlemmarna om pengar . 
De har knappt råd att investera i industrin , än mindre i politiska medel . 
Var inte så självbelåten . 
Hitta sätt att skaffa mer pengar . 
Seongmin . 
Hur många aktier äger du i Seohae Olja ? 
Runt 30 procent , herrn . 
Kan du ge dem till mig ? 
Ursäkta ? 
Jag gör det värt besväret sen . 
Men ändå ... Mina aktier är för ... 
Du kom med i Nationalförsamlingen . Det är ett lågt pris . 
Du behöver mig väl ? 
- Hörde du allt ? 
- Ja . 
Hur många aktier äger du i Seohae Olja ? 
Jag äger 32 procent . 
Vet du vad ? 
Med 62 procent kan du gå med i Cheongwooförbundet . 
Det vågar jag inte . 
Jag ger dig mina aktier . 
På ett villkor . 
Skaffa alla politiska medel . Och i gengäld hjälper jag dig in i Cheongwooförbundet . 
Segangs Textilier Ceremoni för hamnutveckling År 1957 Busan , Sydkorea 
Hej , jag är ledamot An Minchul . 
Min dröm är att sätta Korea på exportkartan . 
Även president Rhee är intresserad av vårt hamnutvecklingsprojekt . 
När hamnen är klar blir Korea ett exportcentrum inom fem till tio år ! 
Uncle Samsik 
Uncle Samsik 
Kallblodig 
Jag var nyfiken på dig , Kim San . 
Jag vill se om du är mer användbar än Kang Seongmin . 
Har du tid att vänta på att bli ledamot och minister ? 
Gör general Choi president så får du makten direkt . 
Håller du inte med ? 
Det är väl det du vill ? 
Vet du att Kang Seongmin dödade min storebror ? 
Farbror Samsik . 
Farbror Samsik . 
An Kichul vet allt . 
Ursäkta ? 
Om vem som dödade An Minchul . 
Vad menar du ? Vet han att det var vi ? 
Han vet allt . 
Förlåt , men jag råkade nämna uppförandekoden . 
Berättade du om uppförandekoden ? 
Du borde träffa An Kichul . 
19 mars 1960 Seoul , Sydkorea 
Hotell Banya 
Utgången är till vänster . 
Jag såg många utlänningar i korridoren . 
Vilka är de ? 
Inspektörer från FN . 
Kom in . 
Tog du med den ? 
Ja . 
Signaturen är tydlig . 
Verkligen . 
Farbror Samsik . 
När hotellet byggdes var det här min fars kontor . 
Jag brukade rusa in och ut hela tiden . 
På den tiden verkade hotellet enormt . Men nu verkar det så litet . 
Det är fortfarande Koreas bästa hotell . 
Precis . 
Korea är för litet för mig . 
Stöttar du familjen An eller familjen Kang ? 
Ursäkta ? 
Givetvis stöttar jag familjen An . 
Skönt att höra . 
För de två familjerna har blivit osams nu . 
Jag förstår . 
Jag visste att Kang Seongmin dödade min bror . 
Din metod funkar inte för utbildade människor . 
Den funkar bara för folk som Yoon Palbong . 
Min far sa alltid att du skulle bli användbar . 
Jag förstår . 
Jag ska göra mitt bästa . 
Hur inblandad var du i mordet på min bror ? 
Jag förde bara Yoon Palbong till Busan . 
Jag trodde aldrig att Kang Seongmin skulle mörda ledamot An . 
Efter kuppen kommer Kang Seongmin att avrättas lagligt . 
Är du redo för det ? 
Du har en dålig vana . Du underskattar yngre motståndare . 
Du måste ändra på det . 
Det ska jag . 
Tack för ditt vänliga råd . 
Jag menar inte mig själv . 
Jag menar Kim San . 
Underskatta honom inte . 
FN-inspektörerna är här . 
Vad sa An Kichul ? 
Kolla upp An Kichul . Vi måste krossa honom . 
Vad är det nu ? 
Vi kan inte låta honom vara . Doochill . 
Glöm det . Tiderna har förändrats . 
Våra metoder funkar inte . 
Varför har du blivit så svag ? 
Vet du inte vem jag är ? 
Vi måste krossa An Kichul , okej ? 
Jag har känt An Kichul sen han var en bebis , men jag kände honom tydligen inte alls . 
Jag visste inte att han var listigare än sin far . 
Den pojken är inte lika bra som sina äldre bröder . 
Han är fortfarande ung och ödmjuk . 
Ni måste ta hand om honom . 
Inte ens hans egen far genomskådade honom . 
Kan vi lita helt på Kang Seongmin ? 
Nej . 
Inte ? Har du några idéer ? 
Ja . 
Jag har en storslagen plan för hur Cheongwooförbundet ska ta över landet . 
En storslagen plan ? 
Vi inför ett parlamentariskt system och mutar hela Nationalförsamlingen . 
När jag presenterade min plan måste snorungen ha skrattat åt mig . 
Kan du gå ut ? 
Det var väl meningslöst eftersom jag inte kunde avvisa Kang Seongmin . 
Minchul uppnådde inte sin dröm . Låt mig förverkliga den . 
Jag kan göra det . 
Svär du på att du inte dödade min son ? 
Han såg nog ner på både Kang Seongmin och mig . 
Vem dödade då min son och varför ? 
Jag ska ta reda på det . 
Jag ska gå till botten med det . 
Herrn . 
Om Cheongwooförbundet överger mig har jag ingenstans att ta vägen . 
För att han har sett oss kräla vid hans fars fötter . 
Jag ska vara lojal . 
Snälla , hjälp mig den här gången . 
Bara den här gången . Skona mig . 
Hur ska du bevisa det ? 
Jag gör vad som helst . 
- Vad som helst ? 
- Ja , vad som helst ! 
Om jag bara hade sett hans blick ... 
Hur kunde jag missa det ? 
Missa att An Kichul var kallblodigare än Kang Seongmin ? 
Utvecklingsbanken beviljar oss ett lån för lokalerna , varav 30 % kommer att användas till valkampanjen . 
Va ? 30 % ? 
- Det är absurt . 
- Otroligt . 
Det är för mycket . 
När jag tar över valkampanjen ska Liberala partiet ledas av Cheongwooförbundet . 
När det händer kan vi yrka på en lag gällande industrikomplexet . 
Lita på mig och visa ert stöd . 
En applåd ! 
Han måste ha hånat oss inombords medan han iakttog oss i tysthet . 
Alla drömmer om absolut makt . Men saken är den att om nån kan reformera politiken varför inte bli president ? 
Kim San hade inte en chans mot den sluga lilla ormen . 
Gör general Choi president så får du makten direkt . 
Sn Kichul kan vara oemotståndligt lockande . 
Det är väl det du vill ? 
Kim San är ingen match för honom . 
Du är mycket bättre än Kang Seongmin . 
Men An Kichul skulle ha insett Kim Sans värde . 
Farbror Samsik vill göra Kang Seongmin till premiärminister . 
Kan vi införa parlamentsystemet ? 
Jag vet inte . 
Jag tvivlar på det . 
Det sa jag till min far också . 
Det är Kim Sans svaghet . 
Så varför ... 
Det var vad min far ville . 
Men inte vad jag vill . 
Kim San dras till folk som inser hans värde . 
Varför ville du träffa mig ? 
Jag var nyfiken på dig . 
Jag vill se om du är mer användbar än Kang Seongmin . 
Varför gör du dig sånt besvär ? 
Döda mig direkt . 
Det vill jag gärna . 
Försöker An Kichul rädda Kim San ? 
Han gjorde en begäran till revolutionsarmén . 
Så du lyckades övertala general Choi ? 
Det stämmer . 
Varför ändrade han sig ? 
Han ändrade sig inte . Jag ändrade mig . 
Ministeriet för rekonstruktion då ? 
Blir det inget ? 
Jag vill etablera det . 
Jag tänker göra det själv . 
Jag struntar i parlamenssystemet och kuppen . 
Och jag trodde aldrig på politikerna . 
Han ser bekant ut . 
Kim San struntar i vem som tar makten så länge han kan realisera rekonstruktionsprojektet . 
Demokraterna är splittrade mellan Yoon Bohyuns gamla och Jang Mins nya grupp . 
Jag känner till det . 
Jag vill att policyn hanteras av den nya gruppen . 
Det är enda sättet att vinna den nya partigruppens fulla stöd . 
Dags att rösta om ändringen av lokalt självstyre . 
Att hyllas som demokratins väktare ? 
Kom igen . 
Det var Kim San aldrig intresserad av . 
- Hur vågar ni ? - Vi knuffar oss in . 
Håll armkrok ! 
Lagförslaget är ogiltigt ! 
Inga illegala val ! 
- Lagförslaget är ogiltigt ! 
- Vad i ... Släpp . 
Inga illegala val , Kang Seongmin . 
Hur vågar du attackera en ledamot ? 
Du är ingen ledamot . Du är Choi Minkyus lakej . Din lilla ... 
- Herrn . - Vi fördömer starkt att lagförslaget antogs så skyndsamt och begär en officiell ursäkt till ordförande Kim San . 
Det skiljer Kim San från Kang Seongmin . 
Det är onödigt . 
Jag godtar hans ursäkt . 
Va ? 
- Du kan inte släta över saker . 
- Jo , ibland . 
Det räcker . 
Den 3 april 1960 Seoul , Sydkorea 
FN-inspektörerna ska utreda valet . 
De föreslår nog en omröstning . 
Har det nåt inflytande ? 
Det sätter press . 
Du kan väl vänta lite till ? 
Du kan uppnå ditt mål även utan en statskupp . 
All väntan kommer att kosta dig din chans . 
Statskuppen kommer att omvälva koreansk politik . 
Vi behöver ett rättfärdigande . 
En revolution kräver mer än beslutsamhet . 
Kliv in . 
Hej . 
Jag är kapten Lee Sooil från 55:e Howitzerregementet . 
Kapten Lee Sooil från 55:e Howitzerregementet ? 
Tack för att du kom . 
Överste Baek Hyunseok från underrättelsedivisionen ? 
Jag är överstelöjtnant Jeong Hanmin . 
Tack för att du kom . 
Var är general Choi ? 
Han är på en säker plats . 
Är det på hans order ? 
Jag följer hans direkta order . 
Kliv in . 
11 april 1960 Masan , Sydkorea 
Masans kust 
Daegus studentprotester är våldsamma . 
- Nåt nytt om Masan ? - Inte än . 
Jag är Cha Taemin . 
Nån stal valurnorna där oppositionen ledde . Men vi hittade dem . 
Och jag vill be om ursäkt . 
Yoon Palbong , Kim Kwangmin och Kim San . 
Nån står bakom dem . Nån utmålade min far som ett monster . Nån fick bort mig från säkerhetsbyrån . 
Nån fick min far dödad , anklagade honom för att vara spion och gör San till ett monster . 
Far . Bjöd du in liberala ledamoten Pak Jiwook ? 
Han ringde tidigare . 
Men han torterade dig under den japanska ockupationen . 
Du har rätt . 
Men nu är jag politiker och måste släppa det . 
Jag vet inte var jag ska börja , men Pak Jiwook satte dit flera oskyldiga medborgare under japanskt styre . 
Vem var bakom Yoon Palbong ? 
Det kan jag tyvärr inte berätta . 
Så du vet . 
Enligt polisrapporten sköts Yoon Palbong först . 
Även andra skottet var riktat mot honom . 
Vad betyder det ? 
Ska vi bara låta det vara med alla obesvarade frågor ? 
Det är farbror Samsik , va ? 
Stal ni valurnorna ? 
Inget om Masan ? 
Nåt från herr Kim ? 
Det är min son ! 
Låt mig se honom ! 
Min stackars älskling ... 
Vad hände ? 
Min stackars älskling ! 
Såg du kroppen ? 
Ja , han kastades i havet med en tårbomb i ansiktet . 
Va ? 
Aemin Dagblads politikavdelning . 
Vem är det som ringer ? 
Yeojin , det är till dig . 
- Vem är det ? 
- Jag vet inte . 
Choo Yeojin . 
Jag är Cha Taemin . 
Jag tror att Pak Jiwooks män är där borta . 
- Håll dem borta . 
Ursäkta mig . 
- Hej . 
- Ursäkta mig . 
Vart är du på väg ? 
- Släpp fram mig . - Vänta . 
Du är bekant . 
Släng allt som har med valet att göra ! 
Det finns inget att tänka på ! 
Kasta allt som rör valet ! 
Är ni osäkra ? Tänk inte och ställ inga frågor . 
Bara bränn allt ! 
Fortsätt så , nu kör vi ! 
Den här vägen . 
Tack för att ni väntade . 
FN-inspektörerna kommer i morgon . 
Svara på deras frågor . 
Upprepa att du inte vet nåt . 
Hur kan du vara så lugn ? 
Vi är körda om de inser att vi stal valurnorna . 
Gör dig av med Samsik . 
Va ? 
Att stjäla valurnorna var inte min idé . 
Du drev mig till att göra det och nu ska jag ta konsekvenserna ? 
Vad fan sa du ? 
Din lilla ... 
Stanna där ... 
Den jäveln . 
Det är jag . 
Ser du lastbilen ? 
Valurnorna står i den . Angående din fars incident ... Det var en olycka . 
Jag vet . 
Jag ber om ursäkt . 
Farbror Samsik . 
Hur är han ? 
Han har utnyttjat dig hela ditt liv . 
Jag står för det jag har gjort och hedrar alliansens kodex . 
Bageri Sail 
Valurna för presidentvalet Cheonjuns vallokal 
Det är jag . 
Journalister går in på Aemin Dagblad . 
Ska jag ingripa ? 
Nej , gör inte det . Avvakta bara . 
De var här ganska länge . 
Överstelöjtnant Jeong Hanmin ? 
Ja , han har varit här förut . 
Titta här . 
Reservationen gjordes av kapitalförsvaret . 
Hur många var de ? 
Runt tio stycken . 
Hörde du vad de sa ? 
Jag hörde en viss general nämnas flera gånger . 
General Choi Hanrim ? 
Ja , det var han . 
Vet du vem mer som var här ? 
Kapten Lee Sooil från Howitzerregementet . Och en överste från arméhögkvarteret . 
Kolla upp kapten Lee Sooil . 
Ja , herrn . 
Herrn . 
Vad är det ? 
Vår position är röjd . Det är farligt att stanna . 
Vi går till bunkern . 
Vem fick reda på platsen ? 
Det måste hamna på förstasidorna imorgon . 
Låt alla journalister turas om att bevaka valurnorna . 
Översätt det till engelska så fort som möjligt . 
Det är bevis på gruppröstning och mobilisering av regeringsarbetare . 
Vi bombarderas med tips . Ska jag summera dem ? 
Inkludera alla bevis på det liberala partiets valfusk i rapporten . 
Det 55:e Howitzerregementet , arméhögkvarteret och 3:e marinkårsregementet . 
Det var nog de officerarna som planerade statskuppen . 
Vad sa Choi Hanrim ? 
Att vi ska vänta på FN:s inspektion . 
Det finns två möjligheter . 
Choi Hanrim har ändrat sig eller ... Hanmin utnyttjar general Choi . 
Det stämmer . 
Vi ses på bageriet sen . 
General Choi är i bunkern . 
Har han bestämt sig ? Ja , herrn . 
Är han inne ? 
Herrn . 
Hallå där . 
Är du knäpp ? 
Ska du be om ursäkt ? 
Be om ursäkt ? Varför då ? 
Lugna dig , herrn . 
Hur kan jag lugna mig om det blir omval ? 
Du kan gå . 
Har du kollat valurnorna ? 
Varför har du inte gjort det själv ? 
Gå och kolla med Samsik . 
Visst . 
Vi måste göra oss av med honom . 
Är det för mycket för dig ? 
Du kan lita på honom . 
Han vet allt ! 
Sluta gnälla , för fan . 
Jag hanterar farbror Samsik som jag vill . 
Säg inte åt mig vad jag ska göra . 
Du är ansvarig för den här röran . Sluta gnälla , så ses vi imorgon . 
Var är general Choi ? Han är där inne . Kom . 
Kapten Lee Sooil på 55:e Howitzerregementet . 
Hans far är vd för Samjin Textilier . 
Samjin Textilier ? Ett dotterbolag till An Yosubs företag . 
Kapten Lee Sooil Han gick på Militärakademin . 
An Kichul måste ha diskuterat kuppen med honom från början . 
Nåt nytt om general Choi ? 
Pak borde vara tillbaka nu . 
Är han inte där ? 
Blev han bortförd ? 
Han blev bortförd . 
Okej . 
Det var nog Hanmin . 
Jeong Hanmins trupper är inte fler än 2 000-3 000 . 
Vad gör vi om USA:s armé ingriper ? 
De är många fler än vi . 
Ja . Tack . 
General Choi är här . 
Tänk om Choi Hanrim fortfarande tvekar ? 
Vi går vidare . 
Jag ska hindra USA:s inblandning . 
- Jag räknar med dig . 
- Okej . 
Hanmin kan inte ha gjort det ensam . 
Kan An Kichul ha övertalat honom ? 
Vad sa An Kichul ? 
Att han skulle döda Kang Seongmin . 
Döda honom lagligt . 
- Med alliansens uppförandekod ? - Ja . 
I den här takten är general Choi i fara . 
Varför ? 
Han föreslog att vi väntar på FN:s inspektion . Men det går de inte med på . 
Om vi inte stoppar An Kichul nu dödar han mig först . 
Han nöjer sig inte med dig . 
Han dödar alla , inklusive mig och Kang Seongmin . 
Efter statskuppen ... 
Herrn . 
Du sa inte att du skulle komma . 
Så nån vill se mig död ? 
Och nåt om en kupp ? 
An Kichul vet allt . 
- Vad ? 
- Att du dödade hans storebror . 
Han vet allt . 
Visste An Yosub det ? Ja . 
Han visste allt . 
Vad menar han med att döda mig lagligt ? 
- Med uppförandekoden ... - Det är inte det . 
Alliansens uppförandekod ? 
Vi brände den . 
Pak Jiwook gömde originalet . 
Pak Jiwook gömde originalet ? 
Ja , herrn . 
Jag varnade dig för honom . 
Han jobbade för japanska polisen . 
Jag bad dig akta dig . 
Valurnorna , då ? 
Tog ni hand om dem ? 
Valurnorna ... 
Saken är den ... 
Cha Taemin tog dem . 
Varför då ? 
För att tipsa Aemin Dagblad , vilket är gjort . 
Ni klantade er med Pak Jiwook och valurnorna och gjorde ingenting när An Kichul försökte döda mig ? 
Förlåt , herrn . 
Vad händer med mig om det blir känt ? 
Jag kan inget säga . 
Du skulle övervaka An Yosub . 
Vad fan har du gjort ? 
Skyll inte på farbror Samsik . 
- Va ? 
- Det är ditt fel , inte hans . 
Han är lite burdus . Förlåt honom . 
Jag säger sanningen . 
Albrightstipendium ? 
Bäst i klassen ? 
Åt helvete med det . 
Vad sa du ? 
Sluta spela oskyldig . 
Du ville krossa mig och ta min plats . 
Trodde du att jag inte visste ? 
Du visste att valurnorna skulle stjälas . 
Varför gjorde du inget ? 
Din jävla hycklare . 
- Du är precis som jag . 
- Jag är inte som du . 
Jag jobbade hårt , vann ett stipendium och allt . 
Mina föräldrar har inte förrått sitt land . 
- Vem hade det lätt ? - Sluta nu . - Ni vet bättre . - Berätta om jag hade det lätt . 
Du vet hur mitt liv var . 
Jag vet mycket väl . 
Vår kära herr Kang har gått igenom mycket . 
Du kan inte undsätta honom jämt . 
Undsätta ? 
Hördu . 
Vem tror du fick farbror Samsik dit han är nu ? 
Det var familjen Kang . 
Du har varit deras slav . 
Han är ingen slav . 
En slav är nån som du . 
Du tror att farbror Samsik ska göra dig fri ... 
Vi har inte tid med detta . 
Vi måste stoppa An Kichul ! 
Bäst att du har en plan . 
Jag har en plan . 
Vad är det ? 
Undantagstillstånd . 
För att förhindra truppförflyttning . 
Det var enda sättet att förhindra kuppen . 
Demokrati stulen ihop med valurnor 
Det var enkelt . 
Aemin Dagblad rapporterade om stölden av valurnorna . 
- Vad i ... 
- Vad hände sen ? 
Helvetet bröt lös . 
Herr president , förklara undantagstillstånd . 
Det råder undantagstillstånd . 
Herrn . 
Det finns ingen återvändo nu . 
Detta är kapitalförsvarets största operation sen kriget . 
Det här är ingen övning . 
Vårt land är en enda röra . 
Vi soldater måste agera . 
Vi ska visa vad vi kan . 
Ingen kommer till skada om vi håller oss till planen . 
Undantagstillstånd ? 
Vems idé var det ? 
Det var min idé . 
