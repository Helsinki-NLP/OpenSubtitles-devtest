Är vi nästan framme ? 
Jag ... Jag har blöta strumpor . 
Det måste vara minus 50 . 
Pappa ? 
Vad ska vi göra nu ? 
Varm choklad ? 
Var ska vi bo , menar jag . 
Tja , vi kan åka hem till England . 
Vi kan stanna här i Sverige . 
Vi kan åka vartsomhelst . 
Jag menar , vi har inga ... Minns du senast vi var här ? 
Det var sista sommaren med mamma . 
Jag är nervös . 
Hon kommer inte att vara här . Det vet du väl ? 
Vi kommer inte att se henne igen . 
God jul i efterskott och grattis på födelsedagen i efterskott ! 
Okej . " Vad står mitt i elden utan att bränna sig ? " 
" Bokstaven D. " 
Den var rätt bra . 
Vad ? 
Den var usel . 
De ska vara usla . Det är poängen . 
Din tur Åh , nej . 
- Jo . - Jo . Din tur . 
Okej . Okej , jag har en . 
Den är lite lik den andra . 
- Men lite svensk . - Jag är gift med en svensk . Varsågod . 
Okej , så , Nelson Mandela har en svensk halvbror . 
Vem är Nelson Mandela ? 
Det funkar inte om du inte vet vem Nelson Mandela är . 
Jag vet vem han var . 
Okej , så Nelson Mandela har en svensk halvbror som heter MåsteMandela . 
Den är jättekul på svenska . 
Du har ändrat om i skåpen . 
Nej , jag är inte direkt typen som ändrar om i skåp . 
Jo , kan vi prata ? 
Självklart . 
Det är bara ... Vår relation var inte direkt den bästa när du åkte . 
Hur var vår relation ? 
Du ... tittade inte på mig ... när vi sa adjö . 
Såklart jag gjorde . Nej . Det gjorde du inte . 
Jag har tänkt mycket på det det senaste året . 
Jag vet inte om du märkte det , men det var några verkligt förfärliga månader . 
För mig , åtminstone . Innan du åkte . 
Jag är ledsen . 
Det är inte så jag minns det . 
Jag är tillbaka för att stanna . 
Älskar du mig ? 
Såklart jag gör . 
Jag är inte bara ömhetstörstande . Det är en genuin fråga . 
Såklart jag älskar dig , din stora idiot . 
- Hej . 
- Välkommen tillbaka , ma ' am . 
Tack . 
Den här , då ? " Hur sanden kom till havet . " 
Slänga eller behålla ? 
Du förstår mig inte alls , va ? 
Jag frågade om du ville behålla eller kasta den . 
Kasta . 
Kastad . 
The Changeling . 
Ja . Den där trollen tar bebisen . 
Och de kastar barnet i elden för att få tillbaka mamman . 
Var det nåt särskilt som upprörde dig innan jag åkte ? 
Vi behöver inte prata om det . 
Har du sett insexnyckeln ? Ja . 
- Det är väl den här ? - Ja . 
Vi såg dig knappt . 
Visst , vi hade den där bortregnade sommaren uppe i stugan , men du var iväg på träning . Mycket . Så det var inget specifikt ? 
Vet du , det kommer en dag då jag har monterat ihop min sista skitmöbel och aldrig behöver göra det här igen . 
Magnus , vad ? 
Jag är ingen svartsjuk person . Det hoppas jag att du vet . 
Men jag hade verkligen börjat undra över dig och Frederic . 
Vad ? 
Absolut inte . Nej . Du , det går riktigt bra mellan oss . 
- Ja . - Så nu vore en bra tid att vara ärlig mot mig . 
Men Magnus , jag var inte otrogen med Frederic . 
Jag skulle aldrig göra så . 
- Visst . 
- Magnus , snälla . 
Jag vill bara att vi är ärliga . Ja . 
Jo , medan du var borta träffade jag nån . 
Vad ? 
Inget hände egentligen . 
Vi gick ut på en drink . 
En kyss . Vad ? 
Jag trodde att du skulle lämna mig , Jo . 
Du vet , det pågick mycket skvaller om dig och Frederic . 
Jag antog att det var slut mellan oss . Men varför ? 
- Alltså ... - Jag försöker bara vara ärlig . Ja . Jag vill att du ska vara min man , okej ? Jag vill att Alice ska vara min dotter . 
Det enda jag kunde fokusera på där uppe var att ta mig hem och montera ihop billiga möbler . 
När jag var där uppe , helt ensam , och ingen kunde höra mig , och jag trodde att jag skulle dö . 
Pappa ? Pappa . Kom . 
Magnus ... Jag sörjer tiden som jag har förlorat med dig och henne . 
Jag skulle inte stå ut med ... Pappa ? 
Förlåt . 
Mr Rogers ? 
- Mr Rogers ? - Ett ögonblick . 
- Är han ... 
- Bud , alla talare ska gå till huvudsalongen för krisinformation . Ja , jag ville bara säga ... Lystring , tack . Mina damer och herrar , det här är kapten som talar . 
Vi ska vända och göra ett stopp i Santa Barbara . 
Det verkar ha skett en incident med en av våra gäster under natten . 
Det krävs några nödvändiga säkerhetsåtgärder och förfaranden . 
Vi ber er stanna ombord , och hoppas att detta inte är en alltför stor olägenhet . 
Henry , du är finansierad och anställd av NASA . 
Och har varit det sen långt innan du föddes , Michaela . 
Vi måste prata om det faktum att du inte fått tillstånd att ta med RPL-utrustning till en annan rymdbyrå . 
CAL är min . 
- Den fungerade inte , Henry . 
- Nej , snälla säg inte så . 
Jag vet . Det är väldigt svårt att släppa taget . 
Det här är inget misslyckande . Jag behöver bara tänka igenom det . Det har en inverkan . 
Du måste komma hem , okej ? 
Du har fått tio dagar med mycket assistans och det finns inga bevis för att CAL funkade . Vi lägger ner . 
Projektet är avslutat . Henry ... Jag minns saker fel . 
Såsom ? 
Var saker finns . Min bil . 
Jag minns den som röd , men den är blå . 
Det är en småsak , men ... Det är faktiskt en ganska stor sak . 
Jag tror att jag ... Jag har ett piano hemma , och jag spelar inte piano . 
Får du hallucinationer ? 
Av vilket slag ? 
Jag ser Paul Lancaster . 
Jag menar , jag ... Hans vålnad , antar jag . 
Ibland känns det som om jag fortfarande är kvar där uppe på ISS . 
Det du har berättat verkar högst symptomatiskt för PTSD , där man skulle vänta sig upprepningar av stressande händelser , minnesluckor , vrede . 
Det vore inte förvånande om du har det . Du fruktade för ditt liv och var väldigt orolig för din besättning , din familj . Hanterade en väns dödsfall . Du har genomlidit ett oerhört trauma . 
Nu är du tillbaka på jorden och börjar känna av effekterna . 
Vi gör ett dexametasonhämningstest för att kolla dina kortisolnivåer . 
Och under tiden kan jag ge dig nåt . Såsom ? 
Litium . 
Jenny , jag är inte psykotisk . Jag är inte deprimerad . 
Nej , men det lugnar ner dig . 
Det lugnar ner såna här saker . 
Jag vill inte det här . Jag är inte ... Sånt här är karriärsavslutande . 
Jag är intresserad av din forskning . 
Vad kallas det , " salutogenes " ? 
- Jag ... - Hur definierar du det ? 
Jag visste inte att du var här . Jo , jag är här . 
Det är nog en bättre plats för mig . Jag tror att jag kan hjälpa . 
Så hur går det för dig ? 
Med CAL , menar du ? 
Jag kör den om och om igen . 
Jag tror att jag kan vara nära ett genombrott . 
Jag minns inte mycket om CAL före olyckan . Jag ... - Jag ... - Vill du se det ? 
Jag får inte in mycket jag förstår . 
Har du hört mycket anekdotisk bevisföring från astronauter ? Hur de påverkas ? Det är inte enbart bra . 
Jag vet att några kände sig utbrända . Ja . 
Folk tycker att det är tufft . 
Upplever saker de inte förstår . Ja . 
Jag har ett par vänner , besättning på Gemini IV , Chuck Parks och John Cooper ... De kände doften av bränt rostat bröd där uppe . Båda två . 
John hörde en hund skälla . 
Sa alltid att det var Lajka . 
Vet du , jag undrar hur Lajka kände . 
Är du hundmänniska ? 
Det har alltid varit fallet sen vi började flyga på höga altituder . 
Jag var testpilot , före Apollo . 
Flög till de högsta möjliga altituderna , ända upp till rymdkanten . 
Det var ganska vanligt på den tiden att kollegor rapporterade en stark kraft som pressade ner en av planets vingar ovanför 27 000 meter . 
De kallade det " Guds vänstra hand " . 
Jag kände en kille . Han hade mist sin son . 
En liten pojke , sex år gammal , som drunknat i en sjö på sin lillasysters födelsedag . 
Några år senare flög killen DC-10:or över Nevada och hörde en röst . 
Sin sons röst . " Pappa , se upp . " 
Han insåg att han börjat störtdyka och lyckades räta upp planet . 
Fram till sin död svor han på att hans son räddade honom . 
De säger det inte , men det är såna saker som följde oss upp i rymden . 
SALJUT 7-BESÄTTNINGEN SOM SÅG ÄNGLAR Har du nånsin sett nåt som inte fanns där ? 
Rymdresor är som att bestiga Everest . All fokus läggs på att nå toppen och om man inte passar sig , kan man glömma att man måste ta sig ner igen när man nått den . 
Det är då folk rasar . 
Jag måste kolla det här . Den är igång igen . 
- Hej . - Det är pappa . Jag kan inte prata . 
Det funkar inte . 
Åh , gud . Det gick bra i några år , men ... Herregud , jag måste hitta en lösning . Jag måste hitta ett sätt att sätta dit den jäveln . 
Du måste sluta tänka som om allt det här finns utanför dig . 
Connie , det är ingen sjukdom . 
Det är en sjukdom . Ingen har mixtrat med din hjärna . 
Det är du . Det är nåt du kan kontrollera . 
Om du har en episod , snälla , ta bara din medicin . 
Som sagt , jag kan inte prata . 
Hon pratar om död och olyckor . 
- Och vi har ett skåpproblem . - Vad menar du ? 
- Hon gömmer sig i skåp . Ja . - Hon gömmer sig i skåp . 
Det verkar för mig som om ni kanske har förlorat varandra lite . 
Hon är tio . Hon var nio när du åkte . 
Det är ett långt år . Det är en väldigt liminal ålder . 
Vad menar du med " liminal " ? 
Mellan en sak och en annan . Ja . Exakt . 
Hon vill ändra om saker , som sitt rum . 
Och i ett år har ni haft fadern och dottern , så mamma är ... Mamma har varit för långt borta . Hon var i rymden . Nu är hon tillbaka , och kanske är Alice inte säker . 
Hon kanske plågas av känslor som : " Mamma är ... Vem är du ? 
Kan jag lita på dig ? " 
Vad har du sagt till henne ? 
Hon känner till privata saker . 
Hon är min kollega och Alices lärare . 
Vad sa Jenny ? 
Jenny sa att jag har PTSD . 
Det är inget att oroa sig för . Jag mår bra . Berätta inte för nån . 
Tror du att det är nåt fel på min anknytning till Alice ? 
- Nej ? Självklart är det det . 
Jag har varit borta i ett år . 
" Vem är du ? 
Kan jag lita på dig ? " 
- Hon sa inte att hon inte litar på dig . 
- Du satt bara där och höll med . 
Kolla i gästrummet . 
Är du här ? 
Alice , kom ut därifrån . 
Alice , nu . 
Vad ? 
Jag har lite gamla kläder som du kanske skulle gilla . 
Älskling . Kom . 
Vi har inte riktigt haft tillräckligt med mamma-Alice-tid . 
Vi kanske kan åka bort nånstans . 
Bara vi två ? 
Nej . Pappa också , såklart . 
Vi kan åka till stugan . 
Men skolan , då ? 
Skolan har haft dig i ett helt år . 
Älskling , stäng inte mig ute . Det gör jag inte . 
Är du inte glad att jag är hemma ? 
Jag vet inte . 
Jag är bara lite besviken . 
Jag trodde det skulle bli annorlunda . 
Mitt i CAL finns en kammare innehållande en gas av rubidiumatomer . Runt den finns lasrar , elektromagneter . 
- En magnetisk fälla . - Förstått . För att få kondensatet riktas lasern för att ge resonans av atomerna . 
Sen , när lasern stängs av , det är då överlagringen bildas . 
Bildade ni den ? 
En svart konturlös massa ... Två svarta massor jämsides . 
Det här är bilden vi fick ombord på ISS . 
Det finns en interferenseffekt , Henry . Det får inte finnas en interferenseffekt . 
Vad visar uppgifterna nu ? 
- Här . - Vad är det här ? Det ser ut som en barnteckning av en uggla eller nåt . 
Det vill inte bli sett . Vad ? 
Men tro mig , när jag har haft igång den här nere ... Haft igång den här nere ? Så är det vad jag ser . 
Visa mig uppgifterna då . 
Det här är uppgifterna . Jag kan inte , Louis . 
Det finns där , klart och tydligt , inuti glorian , men bara jag kan se det . 
Ledsen , Henry . Du kan inte ha byggt en portal till ett annat universum . 
Det du såg från ISS var en falsk bild . Nej . CAL-experimentet var ämnat att fånga ett tillstånd i vilket en partikel befinner sig i två olika tillstånd samtidigt . 
Och vi gjorde det . 
Henry , ett experiment gick snett och du fick en falsk bild . Men du kan alltid försöka igen . 
Nej , sir , Jag kan fanimej inte försöka igen , för vi kommer aldrig att åka dit igen . 
Lyssna , Louis , tänk om resultatet av experimentet teoretiskt kunde synliggöra sig på olika sätt . 
Såsom ? 
Inte på en skärm . I sinnet på en observatör . 
Av vad du ser i världen runtom dig . Tänk om det påverkar hjärnans kemi ? 
Snälla du . Hela kvantumfysikens historia är nära förbunden med observatörseffekten , hur experimentet påverkas av att nån tittar på nåt . 
Tänk om experimentet påverkar mig ? 
Det måste väl göra ont ? När nån inte tror er . 
Agent Bright , FBI . 
Ni vet att det vi diskuterar här är en psykologisk sjukdom där personerna inte kan se verkligheten som den är . 
Det kan ha undgått er , agent Bright , men sanningen är en bristvara . 
Har det undgått er i rättsväsendet ? Nej . 
Jag var på månen . Jag gick där . 
Det finns bevis . Jag lämnade en golfboll . 
Ingen betvivlar att ni gick på månen . 
Vi vill bara veta vad som hände mannen på fartyget . 
Ni kom och avbröt hans middag . 
För att prata med honom . Få honom att komma till sans . 
De ska släppa av mig i Santa Barbara , okej ? 
Ni sa nåt i stil med att om mr Rogers bråkade med er , så skulle ni kasta honom i havet . 
Nej , agent Bright , jag har inte kunnat lyfta axeln över 45 grader sen jag kraschade mitt plan i Korea . 
Och även om jag kunde , så skulle jag inte . 
Jag är astronaut . 
Det rätta virket . 
Vad gör du ? 
Jag är en oberoende människa . 
Jag behöver ingens tillstånd för att vara nånstans . 
För helvete , jag vill att vi enas om vad som orsakar det här . 
Övertyga mig om att jag inte håller på att bli galen . 
" Ilja . A-vitaminer . " 
" Audrey . A-vitaminer . " 
" Yaz . A-vitaminer . " 
" B-vitaminer . " 
" Amanda Klein . " 
" B-vitaminer . " 
" NASA-astronaut Amanda Klein såg änglar i rymden . " 
Kom igen . 
" Kanadensisk astronaut inför rätta . 
Antog falsk identitet före mordförsök på ex-make , ny familj . " 
" Caldera , Henry . " 
Vad gör ni ? 
Hörni , sluta ! 
Vad jag gör här med min egen tid och mitt eget liv angår bara mig . 
Ursäkta mig , Henry . 
Om du inte hade varit så jävla nyfiken , hade inget av det här varit ett problem . 
Är du okej , Henry ? 
Befälhavare Caldera ? 
Nyfikenhet dödade katten . 
Vi hade mycket tid att fundera , båda två och ingen tid att prata . 
Om vad ? 
Uppenbarligen har nåt förändrats , och jag är ledsen om jag sa saker som var opassande . 
Men jag vill ha dig , Jo , lika mycket som förut . 
Jag vill att vi uppfyller kontrakten här och startar eget , som vi sa . 
Jag har pratat med dem . StarCosm , Alyanna . 
De gillar idén . Särskilt om det är vi två , som ett paket . 
Kalifornien . 
- Jag vet inte vad du pratar om . 
- Jo , hör på . 
Du är skyldig mig att tala om om du har ändrat dig . 
Har du ändrat dig ? 
Det är många konstiga skillnader mellan jorden och rymden , och det är inte bara tyngdkraften . 
Tiden går olika fort på jorden och i rymden . 
Så efter sex månader i rymden , har en astronaut åldrats 0,007 sekunder mindre än en person på jorden . 
Vad händer med den ? 
- Med vad ? - Vart tar de 0,7 sekunderna vägen ? 
Är det du ? 
Ja , jag pratar med dig . 
Är det hon , Magnus ? 
Vad händer ? 
Är det hon ? 
Snälla , Jo . 
- Jag är ledsen , Sara . - " Åh , jag är ledsen , Sara . " 
- Lämna min man ifred , okej ? 
Vad fan var det där ? 
Ge mig nycklarna . 
Det här är löjligt . 
Du skulle inte köra på ett par veckor . 
Jag vet för fan hur man kör en bil . 
Svär inte framför vår dotter . Du beter dig som stans fyllo . 
Kan vi sätta på en sång ? 
Jag måste bara koncenterar mig lite . 
Jag sa att jag måste koncentera mig . 
Alice , stäng av . Stäng av , Alice ! 
- Alice , för helvete . - Mamma ! 
De olika rymdbyråerna har rehabkliniker för astronauter som ... Det finns ett tillstånd som kallas astronaututbränning . 
Hon kom ju just hem . - Hon kan inte åka iväg igen . 
- Hon har ett problem . 
Det är uppenbarligen en reaktion på stressen av det som hände i rymden . 
Och utan ingripande lär hon bli värre . 
Och ska du följa med henne ? 
Jag vet inte . 
Ja , kanske . Till en början . 
Hade du en affär med henne ? 
- Vad har hon sagt ? - Strunt i vad hon har sagt . Hade du det ? 
- Vad är det här ? 
Du ljög för mig . 
Vad ? 
Han är orolig för att du beter dig på ett ganska ... dissociativt sätt . 
Jag kan tala för mig själv , din skithög . 
Vad har du sagt till honom ? 
Jag berättade sanningen . 
Jag ... Ärligt talat ... jag mindes inte . Jag ... - Hur i helvete glömmer man nåt sånt ? 
- Uppenbarligen har du minnesproblem . Dra åt helvete ! 
Om du har de här symptomen , Jo , kan vi lätt skaffa hjälp åt dig . Jag behöver prata med min man . 
Ut ur mitt hus , för helvete . Stick ! 
Jag är inte galen . 
Frederic , jag jobbar för dig . 
Det här är mitt hem . Du hör inte hemma här . Jag är inte på arbetet . 
Visst . Visst . 
Vi går igenom HR i morgon . 
Men det är skönt att allt det här har dragits fram i ljuset . 
- Jag ljög inte för dig . 
- Jag är ingen jävla idiot . 
Jag mindes inte . 
Jag minns inte . Jag minns inte ! 
Kanske är det här inte samma jävla plats som jag lämnade . 
Den är exakt densamma , Jo ! 
Det är du som är annorlunda . Pappa ! 
Vänta . Magnus ! Du , Magnus ... Varför försöker du inte ta hand om ditt barn som omväxling ? 
" Marinobservatoriet . Danmark . " 
" Bästa befälhavare Ericsson bifogat finner du två bandinspelningar . 
Vi hörde er på ISS 15 oktober . 
Inspelningen är inte tydlig , men vi skickar med en transkribering . " 
Vad fan är det för fel på dig ? 
Det är du som säger att du gick på månen och det gjorde du inte . Du är en lögnare , ynkrygg och tjuv . 
- Videorna från SS Bernice är klara . - Toppen . Det är framspolat . 
" TsUP , Stationen här . Snälla svara . " 
TsUP , Stationen här . Snälla svara . 
TsUP , Stationen . Snälla kom . 
Jag ska prata . Jag ... Vet inte om ni hör , men det lyser här , så jag ... Jag vet inte . Jag vet inte om felen finns här eller ... Pappa ? " ... sista transkribering . " 
" Den andra inspelningen gjordes av oss 23 november 1967 . Den verkar visa en olycka i rymden då en kvinnlig kosmonaut dog . " 
Mamma ? 
- Alice ? Vad är det ? Alice ? - Det är jag ! 
Vad ser du ? 
Du var död . 
- Väck henne inte . - Hon är vaken . 
- Det är Wendys pappa . - Vad ? Paul ? 
Snälla , Jo , låt det bara vara . 
- Jag vill gå . - Kom här . 
- Vänta , nej . Sätt ner henne . - Kom här . Kom . Magnus . Vart tar du henne ? 
Sätt henne inte i skåpet ! 
- Sätt henne inte i det jävla skåpet ! 
- Jag vill det . 
- Hur ska det göra saker bättre ? 
- Jag vill att pappa nattar mig . 
- Lägg henne inte i skåpet , för fan ! 
- Hon är rädd för dig , Jo . Okej ? Du skrämmer henne . 
Försvinn bara . Gå ner . 
Jag menar , vad sysslade du med ? 
Varför lägger du henne i skåpet ? 
Hon är rädd . Hon vill gömma sig . 
Hur länge har hon varit rädd ? Hur länge tror du ? 
Ta tabletterna som Jenny gav dig . 
Vet du vad ? - De där tabletterna är antipsykotika . - Självklart . Det är poängen . 
Nej , vänta . Jag menar , båda är det . 
Vitaminerna och ... Båda två ... Det pågår en gemensam ansträngning för att få mig att ta antipsykotika . 
De vill förneka vad jag såg där uppe . 
Ta för fan bara tabletterna , Jo . 
Vad gör du ? 
Jag ska ringa Frederic igen , för han har faktiskt rätt . 
Nej , jag måste reda ut det här . Och du måste hjälpa mig . 
Jag måste reda ut varför de gör så här . 
Jag hjälper dig , Jo . 
Varför ringer du Frederic ? 
Det var ju jag som påstods knulla honom . 
Låt bli ! 
Jag vet att ni alla kunde höra mig när jag var där uppe . 
När jag var där uppe och försökte ta mig hem och var rädd , kunde ni alla höra mig . Jag har hört banden . Och ni tänkte lämna mig att dö där uppe . Jo . 
- Lägg ner telefonen . - Jag är ledsen . 
Lägg ner den jävla telefonen . - Jag kommer att finnas kvar här ! - Lägg ... 
