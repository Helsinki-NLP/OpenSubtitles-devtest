Mamma , vart är vi på väg ? 
Det finns en annan stuga tvärsöver sjön . Kom . 
Raring , vad gör du ? 
Vi måste fortsätta . 
Jag lämnar spår som Hans och Greta . 
Minns du ? Du brukade läsa Hans och Greta för mig . 
Det finns en annan stuga . Som vår stuga , men den är inte vår . 
Vi kommer inte att gå vilse . Kom . 
Mamma ? Mamma ! 
Hon ser inte ut som sig själv . 
Hon är fortfarande din mamma . 
Hon ser död ut . 
Hördu , Alice . 
Tänk om hon inte kommer ut . 
Jag vill ta ett ögonblick för att minnas vår kollega och vän , befälhavare Paul Lancaster . 
Han var en oerhört fantastisk , rolig , hängiven , smart person , en kärleksfull make och far , en fantastisk ledare . 
Och inga ord kan beskriva hur mycket vi saknar honom . 
Era frågor , tack . 
Vad tror ni personligen orsakade olyckan ? 
Det var en kollision . 
Ja , men med vad ? 
Förmodligen nåt väldigt litet . 
ISS har system som skannar efter rymdskrot . 
Det gick ett larm . Vi hann bara inte ... 
Vi är mitt i en gemensam utredning och vill inte förekomma förhören . 
- Ursäkta avbrottet , Jo . - Ingen fara . 
Är ert uppdrag över ? 
Får ni tillbringa lite tid med familjen ? 
Nej , mitt uppdrag är inte över . 
Jag har nio månader av experiment och datainsamling som jag ... Mitt specifika uppdrag har varit att övervaka de fysiska och neurologiska följderna av långvariga rymdresor och ... 
Och känner ni för närvarande de följderna ? 
Jag känner ... Jag känner mig mycket bättre än för några dagar sen . 
Men ni vet man glömmer hur jorden luktar . 
Det finns inget väder i rymden . Inga årstider . 
Så det är väldigt skönt att känna hösten och doften av regn . 
Jag är väldigt glad över att vara hemma . 
Är ni okej ? 
Toppen . Titta , vi är tre igen . 
- Var ska han begravas ? 
- Jag vet inte , raring . 
NASA : S INKVARTERING STAR CITY , RYSSLAND Arlington ? 
Det är där de begraver personer som Neil Armstrong , president John Kennedy . 
Personer från förr ? 
Människor som kommer från USA som har gjort nåt riktigt modigt och viktigt . 
Hjältar som din pappa . 
Erica , han var en fantastisk man . Jag är så ledsen . Frida är mitt namn . 
STAR CITY LABORATORIER STAR CITY , RYSSLAND Vi tog med maskininlärningsgrejerna , det vi kunde bära . 
Det är inte idealiskt , men ... Det spelar ingen roll . Titta . 
Det här är vad vi såg precis innan kollisionen . 
Det finns en interferenseffekt . 
Jag såg samma sak när jag extraherade våra data här nere i Bajkonur . 
- Vad ? 
- Exakt samma . 
Hur då ? Den fungerar bara i rymden . 
- Okej , visa mig . - Jag registrerade inte det . 
Jag menar , det tonade ut , men det var där . Jag såg det . 
Jag vet att det fanns där på ISS , men det kan omöjligen ha överlevt på jorden . 
- Det är omöjligt . - Exakt , Eryn . 
Just därför ska vi utföra det igen med allt det här . 
Välkomna till Berni-Con IV . SCIENCE FICTION-FESTIVAL 2021 
Hej , Bud . Bud ? - Hej . - Vad är ditt traktamente ? 
Fanimej inte nog . 
Tio dagar på ett fartyg , för att prata med några jävla galningar . 
Och kolla in den här killen . 
Jag har gått på den satans månen och så slutar resan så här . 
Jag tvingas sitta och debattera mot den där skitstöveln . - Hej . - Vill ni ha ett glas vatten ? Jag fick 250 . Tjugo dollar per autograf . 
Och mitt i en rymdtragedi . Det är smaklöst . Det är dålig tajming . Och allt förmodat nonsens som hände med mig och de andra ... Fan också . 
Konventkretsen är mycket bättre än skådespeleri . 
Mycket mer sex , till att börja med . 
Jag är less på att höra det . 
Det är så här det är nu . 
Jag är less på status quo . 
Saker kommer att förändras . 
- Hej . - Här kommer utomjordingarna . - Kan du signera till Sophie Space ... - Ja . 
Vi måste viska . Varför då ? 
För att de gör nåt väldigt pillrigt i CAL . 
- Hej , Alice . - Hej , Paul . 
Din mammas stora dag i dag . 
RPL . CAL-data : 
Kärnsignal grön , magneter inriktade , 25,5 . 
- Uppfattat , fas sex . - Uppfattat . 
- Kärntemperatur . - Jag saknar dig så mycket . 
Jag saknar dig med , mamma . Är du försiktig när du går ut ? 
Alltid . 
Jag finner det märkligt att inget MMOD-larm hörs , för jag minns att jag hörde det tydligt . 
Det är viktigt att veta om kollisionen signalerades . 
Och era kollegor , då ? 
Jag minns det inte . 
Det fanns ingen MMOD-datarapport . Inget larm utlöstes . Jag kollade . 
Jag sov . 
Så inget larm utlöstes . 
NASA:s ansvar . Och NASA:s ekonomiska skyldighet . 
Vad är det där för ljud ? Jag har hört det ljudet . Inte bara en gång , utan flera . 
Radiobrus . 
Alla kanaler öppna . 
Besättning samlas i Sojuz 1 evakueringskapsel . Initiera förevakuering . 
Eld och dimma i Zarja . 
- Stäng ner . 
- Houston , det är en brand mellan oss och Sojuz 1 . 
Låt oss samlas i Rassvet istället . 
- Ericsson . - Andrejev . 
- Brostin . - Suri . 
- Jag är fast . - Ericsson , Brostin , luften är klar . 
Kollisionsobjektet visades som ett hinder på elektroniknoden på trussarna . 
Det är inget känt rymdskrot . 
Visa bilderna från rymdpromenaden . 
Jo , sjukvårdsteamet vårdar Paul . Fortsätt rymdpromenaden . Uppfattat . Håll mig uppdaterad . Vart ska jag nu ? 
Instruera henne att gå till truss . Det är avgörande att de lagar de sekundära livsuppehållande systemen . 
Jo , vi ser inte det du ser . Kolla kameran . 
Förstått . Den lyser rött . Det är nåt fel . Tyvärr . 
Vi förlorade video här . Vi har ingen återgivning av vad som hände härnäst . 
NASA / ESA ansvarar för de yttre kamerorna . 
Det uppstod kollisionsskador . Så vi kan inte dra nån slutsats om kollisionsobjektet . 
Det var en kropp . En människokropp . 
Det var en kvinnokropp iklädd sovjetisk rymddräkt och hjälm . 
Kroppen inuti var uttorkad , mumifierad . 
Jag sträckte mig för att röra den . Den lossnade och fortsatte sin omloppsbana . 
Befälhavaren ni inser väl hur osannolikt det är att en kropp har bevarats i rymden i åtminstone 32 år , åtminstone sen Sovjetunionens fall ? Och att ett sånt objekt kunde ha kolliderat med ISS ? 
Självklart inser jag ... Vi har en notering här i våra återställda utskrifter . 
" 06 : 55 : 48 . Ericsson . 
' Kan ni kolla syrgasen ? ' " Vad var ert skäl för att fråga om syrgasen ? 
Det var inga problem med syrgasen i min rymddräkt . 
Testet visar att jag ... Det var inte min fråga . 
Vad var ert skäl för att be om syrgaskontrollen ? 
Jag var orolig för att jag var hypoxisk . Att ni inte fick nog med syre till er hjärna ? 
- Ja . - För att ? 
För att jag , precis som ni , hade svårt att tro det jag såg . 
Ingen kosmonaut eller astronaut har nånsin rapporterats död eller saknad ovanför Karmanlinjen , stämmer inte det ? - Jo . - Så vad är er förklaring ? 
Jag tycker att vi borde börja titta på rymdskrot . 
Har ni varit med om liknande incidenter ? 
Ursäkta ? 
Kände ni att ni upplevde hypoxi , symptom på syrebrist , vid nåt annat tillfälle under ert uppdrag , före eller efter ? 
Symptom på hypoxi inkluderar minnesförlust förvirring hallucinationer . 
Nej . Det gjorde jag inte . 
Kliv av försiktigt . 
Ni ska ta en tablett dagligen tills vidare . 
Vad är det ? 
Folsyra , D-vitamin och B-12 . 
Inget kondensat , bara residuum . 
Det var där . 
Henry , ge dig . Det kan inte ha levt mer än en miljondels sekund . 
" Henry , ge dig " ? Tror du att jag ser ett spöke ? 
Behandla mig inte som en idiot . 
Behandla inte mig som en assistent då . 
Och hur förklarar du det faktum att när jag extraherade data i går , så var det samma bild som vi såg när experimentet utfördes på ISS ? 
Det är en bugg . 
- Det här är ryskt maskineri . - Nu räcker det . 
Ursäkta att jag var kort mot dig , Eryn , men det var fanimej där , även om det inte är det nu . 
Det finns en interferenseffekt . Det finns en koppling , och vi måste ta reda på vad den är . 
Jag gillar din frisyr . 
Jag fäster inte stor vikt vid mitt hår . 
Ju äldre du blir , desto snyggare blir du . 
Dra på trissor . 
Jag fick nog just en komplimang . 
Jag har saknat dig . 
Jag har saknat dig också , Jo . 
Det kändes lite som om jag höll på att drunkna du vet ? 
Förlåt för att jag utsatte dig för det . Nej , nej , nej , nej . 
Vi var överens om det . Eller hur ? 
Vin . 
Jag glömde vinet . 
Pappa ? 
Vad sägs om mamma ? 
Mamma är hemma . Jag vet inte om du hört det . 
Har hon glömt all sin svenska ? Pappa ? 
Vad är det , stumpan ? 
Ett år innan Apollo 11 fanns över 10 000 registrerade fel i kommandokapseln , inkluderande 500 kritiska fel i de livsuppehållande systemen . 
Branden på Apollo 9 orsakades av ett av dessa . Tre människor dog . 
Man hann inte åtgärda problemen innan Armstrong , Aldrin och Collins åkte iväg . 
Förutom , som ni sa , att det gick ett helt år . 
Tror ni att NASA tillbringade det året med att klia sina hemorrojder ? 
Jag vill påpeka , att vi just har mist nån där uppe . En astronaut . 
En verklig person med en verklig familj ... - Punkt fyra , Van Allen-bältet . - Det finns en elementär standard för mänsklig respekt , sir . 
Vi förlorade just hela Internationella rymdstationen ... Med strålningsnivåerna mellan jorden och månen , och kommandomodulens relativa tunnhet , skulle astronauterna ha fått svår strålningssjuka . Ni hade alla dött av leukemi vid det här laget . 
När man lämnar jordens atmosfär , är utträdeshastigheten cirka 16 000 km i timmen . Man passerar igenom Van Allen-bältet på ett ögonblick . 
Radioaktiva partiklar hinner inte interagera med kroppen . 
Så där . Jag deltog . Jag borde inte det , men jag gjorde det . Jag borde ha kastat er i det satans havet . 
Låt mig fråga er en sak . Tror ni att vi är där uppe , eller tror ni att vi bara spelar teater ? 
Vad säger ni , sir ? 
Tror ni att ISS är en saga ? 
Nej . Jag tror att den existerar . 
Jag var inte på Apollo 11 , så jag vet inte om de åkte till månen . Men jag var på Apollo 18 , och vet att jag fanimej gjorde det . 
Ja . Jag har läst er bok . 
Varsågoda , hörni . Boken finns att köpa vid dörren . 
Den är så full av oriktigheter att den är helt värdelös . 
Ursäkta mig ? 
Den är full av sakfel . Till och med namnet på er första hund . 
- Vem skrev den ? - Jag . 
Tror ni inte jag vet namnet på min första hund ? Jag vet inte . Ni får inte rätt på saker , sir . 
Jag tror att ni har tutats i en historia . Eller har ett väldigt opålitligt minne . 
Jag skulle passa mig noga för att kalla mig lögnare . 
Jag tror att ni kanske var på månen . 
Jag tror att de kanske vid det laget hade löst en del problem . Men en katastrof var nära på Apollo 13 , och på ert uppdrag sex år senare , dog två män . 
Jag tror att ni berättar en historia eller så har ni tutats i en historia som inte stämmer . 
Hej , baby ! 
För guds skull . 
Kom igen . Herrejesus ! 
Nej ! Vart fan tar du vägen ? 
Är du okej ? 
Vet inte . Det känns lite konstigt . 
Vill du prata om det ? 
- Det är okej . - Säkert ? 
Ja , säkert . 
Mina ben är så svullna . 
Uppe i rymden , rusar alla vätskor upp i huvudet , och nu forsar de ner . 
Jag hjälper dig . 
Säkert ? 
Okej . Du måste hålla hårt , okej ? - Ja . - Okej . 
- Gick det bra ? - Ja . Försiktigt . Det gick bra . Jag tror du måste gå och hämta pappa . 
Jag är ledsen . 
- Klarar du dig ? - Ja , då . Hämta bara pappa , okej ? 
- Säkert ? - Ja . 
Här . 
Är du okej ? Du föll . Jag hjälper dig . 
Såja . 
Jag är okej . Det är okej . 
En handske tappad av Ed White på USA:s första rymdpromenad . 
En kamera tappad av Michael Collins nära Gemini 10 . 
En räddningsfilt tappad under STS-88 . 
Och de här soppåsarna , kastade överbord av astronauter från Skylab under perioden - 73 / - 74 . 
Jag tror att en soppåse är en bra kandidat . 
Tror ni att en soppåse orsakade olyckan ? 
Nej , jag tror inte att det var en soppåse . 
En soppåses storlek och form ? 
Hade jag sett en soppåse , så hade jag sagt att det var en soppåse , för guds skull . 
Var snäll och behärska er ton , befälhavaren . 
Det är ingens uppgift här att lita på ert ord . 
... elva , 12 , 13 , 14 , 15 , 16 , 17 , 18 , 19 , 20 ! 
Nu kommer jag , beredd eller inte . 
Vi kopierar inte det , hur mycket vi än skulle vilja . 
Kopierar ? 
Jag kopierade det här . 
Det är en teckning , Henry . 
Man vinner inget Nobelpris med bara en teckning . 
Åh , Eryn , det vet jag . 
Jag har redan vunnit ett Nobelpris . 
Ja . Typ 1981 . 
Kan du inte bara hjälpa mig ? 
Fanstyget har varit mitt livsverk de senaste 35 åren . 
Så , varför ser du det men inte jag ? 
Den jädra observatörseffekten . 
Hittad ! 
Vad gjorde du med min kanin ? Det är min kanin . 
- Jag gjorde inget med din kanin . - Varför är du taskig ? Du kan inte vara ond mot nån annans kanin . 
- Jag har din dumma kanin . - Men varför gjorde du det ? Du kan inte göra vad som helst bara för att din pappa är död . 
Det borde ha varit din mamma . 
Din mamma är en galen satmara . Det är vad min mamma sa . 
Din mamma är också en satmara . 
Titta bara på den här diabilden . 
Det här är en soppåse kastad överbord från Mir av sovjetiska kosmonauter . 
NASA uppskattar att cirka 350 av de här är ... 
Befälhavaren , ingen hyser annat än respekt för er och det ni gjorde . Men sekretessen för hela det sovjetiska rymdprogrammets historia har hävts , och det finns dussintals memoarer från kosmonauter , ingenjörer och flygledare som har vittnat , även efter Sovjetunionens fall . 
Vi vet vilka som ingick i kosmonautteamen , vilka som flög och inte , och när de flög . 
Det finns inte enda saknad man eller kvinna i nåt av dem . 
Ni såg nåt som inte fanns där . 
Ni var enormt stressad . 
Det händer . 
Vi ajournerar för i dag . 
Du , jag sticker ut hakan för dig . 
Det gynnar inte oss om det här avgörs av huruvida du fick nog med syre till hjärnan . 
De kommer att fortsätta försöka få dig att verka opålitlig , för de vill inte erkänna möjligheten att nåt av deras rymdskrot orsakade kollisionen . 
Jag såg vad jag såg , för helvete . 
Tar du dina vitaminer ? 
Vad gör du ? 
Jag vet inte vad fan ditt problem är , Jo . Få bara ordning på din redogörelse . 
Magnus ! 
Jag har dig . 
Jag vet inte vad som pågår . Jag känner mig inte som mig själv längre . Okej , nu ser vi bara till att få in dig . 
- Va ... - Här , sätt dig . Det känns som om de attackerar mig hela tiden . 
- Jag vill bara hem . - Okej . Jag vet . 
Låt oss bara ta det försiktigt . Okej ? 
Vill du ta av dig skorna ? Okej . 
Så där . Okej ? Det var en . 
Jag älskar dig . 
Jag älskar dig också . 
Kan du stå upp ? 
Bara ... Sådär . 
Okej . Är du okej ? 
Lyft armen . Såja . 
Där är du . 
Hur mår du , Alice ? 
Jag vet inte . 
Nåt som tynger dig ? 
Åkte du till månen ? En gång . 1977 . 
Hur var det ? 
Ganska bra . 
Vad gör du här ? 
Forskningsgrejer . Som vadå ? 
Har du hört talas om kvantumfysik ? Ja . Jag vet inte vad det är . 
- Vill du veta ? 
Länge styrdes vår förståelse av världen av vad som kallas klassisk fysik . 
- Vet du vad det är ? 
Det är ett elementärt sätt att mäta och förutspå saker . 
Sen kom personer som Albert Einstein . 
- Har du hört talas om honom ? 
- Ja . Ja . Han började forska i riktigt små saker som atomer , subatomära partiklar , vågformer . 
Och det började verka som om klassisk fysik inte gällde längre , vilket är mystiskt . 
Det är inte förutsägbart på sätt som vi för närvarande förstår . 
Till exempel , samma sak kan befinna sig i två olika tillstånd samtidigt . 
Det kan vara en partikel , till exempel , exakt samma partikel . Det finns en värld i vilken den partikeln är svart och en värld i vilken den partikeln är vit . 
Och det finns liksom en punkt av liminalt utrymme mellan de världarna , där partikeln är svart och vit samtidigt . 
Och de verkar inte vilja bestämma sig för ett tillstånd förrän nån tittar på dem . 
Det är galet . Tja , det är galet . 
Men det är verkligt . 
Jag uppfann en maskin som vi tog upp i rymden , - och jag hoppades få svar på ... - Funkade den ? 
Jag vet inte . 
Jag tror att jag såg nåt men det verkar inte vilja bli sett . 
Som kurragömma . 
Precis som kurragömma . 
Jag är ledsen att jag ... Jag lämnade dig ensam . 
Verkar jag vara densamma , tycker du ? 
Inte riktigt . 
Varför ? 
Du ser lite annorlunda på mig . 
Hur ser jag på dig ? 
Som om du gillar mig . 
- Jag tog hem nåt åt dig . - Nämen hej . 
Och jag vill tacka dig för att du tog hem min baby . 
CAL var inget ESA-experiment . Du behövde inte hjälpa mig . Jag uppskattar det . 
- Jo Ericsson . - Henry Caldera . 
Vi har träffats . Ja . 
Du deltog i ... Apollo-programmet . 
Hela mitt liv . 
CAL , det här experimentet , är det viktigt ? 
Det är det för mig . 
Det är stora byråkratier involverade här , befälhavaren . 
Alla har sina egna agendor . Inte bara ryssarna , alla . 
Det är lätt att hamna i kläm . 
De som faktiskt har varit där uppe , de måste skydda sig själva . 
Om du nånsin vill prata ... Tack . 
- Jag trodde du var hos Wendy . - Vi bråkade . 
- Om vad ? - Hon sa att hennes mamma ... Att hennes mamma tycker du är galen . 
Jag hittade rymddräkten som jag tror att det var . 
Den jag såg . Som kolliderade med oss . 
Titta , den ... Det är en Star City-dräkt från början av 60-talet . Saljut 7 och framåt . 
Vet du vem det där är ? Vem ? KVINNLIG KOSMONAUT ÅTERVÄNDER FRÅN RYMDEN Irena . 
Jag säger inte att det var hon . 
Men om det var ett misslyckat sovjetiskt uppdrag , skulle de ha mörkat det . 
Vet ni , jag hörde av en kille att Gagarin inte var först i rymden . 
Det var ... Nej , verkligen . Det var Vladimir Iljusjin . 
Men han störtade i Kina , så de tog hem honom och fängslade honom . 
Det är en konspirationsteori . Vi kan inte börja med konspirationsteorier . 
Det här är ingen konspirationsteori . Det är vad jag såg . 
Vilken är den minst pålitliga formen av bevis ? Audrey . 
Vilken är den minst pålitliga formen av bevis , Jo ? 
Ögonvittnesmål . 
Du är forskare . Du vet det . 
Här är det . 
Det ser dött ut . 
Det repar sig till våren . 
Här . 
Får jag vara ensam en stund , tack ? 
Visst . Ja . 
Någonstädes i rymden hänger mitt hjärta . 
Gnistor strömma ifrån det till andra måttlösa hjärtan . 
Där har ni en av Mirs soppåsar för medicinskt avfall , som de använde på 1980-talet . 
Det finns fortfarande hundratals i omlopp . 
De är väldigt lika . Vi kan godta det här . 
Sovjetiskt rymdskrot , inte vårt ekonomiska ansvar . 
Man måste ta hänsyn till det oerhörda trauma ni alla upplevde . 
Upprepa det . 
Visst . 
Återkallar du ditt påstående om en rymddräkt ? 
Vi är väldigt glada över att vi har konsensus . 
Toppen , Jo . Bra jobbat . 
Får vi åka hem ? 
Har vi ny bil ? 
Vad ? 
Varför gjorde du så ? 
Jag trodde det skulle sväva . 
Du släppte det på golvet som en total dåre . 
Alice , vill du bära upp din väska ? 
- Mår du bra ? - Ja . 
Har vi ny bil ? 
- Vad ? 
- Den är blå . 
Det är den . 
Den är inte röd ... Jag är rätt säker på att vår bil var röd . Nej , den är blå . 
När är sista gången vi gör det här ? 
Det gör mig märkligt bättre till mods . 
Som du sa . 
Drömmer du om jorden eller rymden ? 
Jag drömmer alltid om rymden . 
Jag drömmer om att ändlöst kretsa runt jorden . 
Undrar du varför det är så ? 
Du döljer nåt , Irena . 
Varför är det så viktigt att det inte fanns en död kosmonaut ? 
För att det inte fanns nån död kosmonaut . 
Kanske fanns det det . 
Jag är döende ... Jag har lymfkörtelcancer . Stadium fyra . 
Så det här är sista gången . 
Är du verkligen döende , Valja ? 
Musik . Du får välja . 
Känner du dig märkligt sämre ? 
Allvarligt ? 
- Sen olyckan ? 
- Självklart känner jag mig sämre . 
Jag vet inte vad som kommer att hända mig . 
Jag är orolig att det inte kommer att finnas nån himmel eller nåt helvete . 
Ursäkta . 
- Vill ni göra oss sällskap ? Jag vill att ni går en sväng med mig . 
Inget annat returflyg hade landat inom 160 mil från den avsedda landningsplatsen , men ni lyckades landa en pilotlös modul på 460 meters avstånd från var USS Franklin Roosevelt väntade på den . 
Ja , jag och två döda kroppar . 
Låt mig fråga er , tror ni att jag dödade dem ? 
Är det vad ni vill ? Utmåla mig som mördare ? 
Självklart inte . 
Men ni svimmade väldigt lägligt under trycksänkningen . 
Säg mig ni hur jävla lägligt det är att vakna upp med liken av sina vänner . 
Vi kommer ingenvart . 
Jag har ett evidensbaserat synsätt . 
- Trettio år som överordnad polisman . - Snälla . Sextio år som militärpilot . - Teoretisk fysiker . Astronaut . - Depressiv . Alkoholist . 
Kan ni hjälpa mig ? Vad ? För ni har rätt . Det finns minnesluckor . Saker jag inte minns . 
- Som vad ? 
- Jag lagade det ... 
Jag lagade allt på Apollo 18 . 
De där killarna levde , och sen plötsligt var de döda . 
Förlåt , hur kan ni ha lagat det ? 
Jag lagade det . 
Vi åkte ända till månjäveln , och jag gjorde inte ett enda misstag . 
- Det var Henrys fel . - Vad ? Femtio år av brandy och tabletter . Henry Caldera . 
- Vill ni hjälpa mig ? - Vill ni backa lite ? För jag borde inte stå här och prata med en otäck jävla skitstövel som ni . 
Vill ni veta hur jag vet att jag var där ? För att jag har ett satans hål i mitt huvud . 
Ni vet inte , för ni genomlevde inte det . 
Inte ni heller . 
- Idiot . - Klåpare . - Nej , nej , nej . - Bedragare . 
Vet ni ... Jag är ingen jävla bedragare ! 
Mamma , jag tror inte att det finns nån annan stuga . 
Jag tror ... Vad ? 
Människor kan se saker ibland när de är upprörda . 
Och människor som har varit i rymden , de har sett saker . 
Jag vill inte såra dig . Jag vill verkligen inte uppröra dig , men jag tror att du har rätt ... 
Jag tror inte att du är min dotter . 
Men om jag inte är det , vem är du då ? 
Vad har du gjort med min mamma ? 
