Han har pistol . 
En amerikan . Han har pistol ... Gå in i huset och ring polisen . 
Fort ! 
Vi vill inte döda dig . 
Vi vill inte döda dig . 
För dig är kriget över . 
När en besättning störtade , försvann de . 
Efter bara fyra månader vid Thorpe Abbotts var 32 av de 35 ursprungliga besättningarna saknade i strid . 
Vi talade inte om såna besättningar . 
Vi som fortsatte att flyga uppdrag efter uppdrag måste gå på tå runt deras minnen . 
En del mannar gick upp i limningen . 
De hade sett för många plan explodera framför dem och för många vänner dö . 
Några drack . Andra slogs . Andra låg runt . 
Om man fick chansen att glömma , tog man den . 
Jag själv ? Jag åkte till Oxford University . 
Bubbles död tog mig hårt , och överste Harding ansåg det lämpligt att jag representerade 100:e vid en konferens mellan de Allierade nationerna . Han anmälde mig , och jag åkte gärna . 
- Har ni nånsin varit i Oxford , kapten ? - Nej . Men roligt att vara här . 
Ni hinner kanske inte se så mycket den här gången . 
Med alla föreläsningar och evenemang som planeras , hinner ni nog knappast lämna campus . 
Det är här borta . 
Det finns representanter för nästan alla allierade nationer och territorier . 
Ni träffar nog en del fascinerande människor . 
Det kom för två dagar sen . Hoppas att det inte är brådskande . 
Min fru . 
Hon kan inte låta en vecka gå utan att skicka ett brev till mig . 
Så omtänksamt . 
Har " sub-altern " A M Wesgate anlänt än ? Min rumskamrat ? 
Inte förrän imorgon , tror jag . Och vi säger " subaltern " . 
- " Subbeltärn . " - Subaltern . 
Okej . Jaha , James , tack för rundvisningen . 
Absolut . God kväll , sir . Ha en trevlig konferens . 
" Subaltern . " 
VÄLKOMMEN TILL COOMBE HOUSE Münster var bara Rosies tredje uppdrag , men det var så hemskt att överste Harding beordrade löjtnant Rosenthal och hans besättning att tillbringa en veckas vila på ett ställe vi kallade " flak house " . 
De har hästar här . 
Kan du rida , Rosie ? 
Judar från Brooklyn rider inte . 
- God morgon . - Damerna . Damen . 
- Hej . - Se upp . Här kommer kavalleriet . 
Välkomna till Coombe House . 
Vi har alla sporter och aktiviteter man kan önska , precis här . 
Vi har tennis , cykling , volleyboll , krocket , rida med hundar . 
Och om det regnar , för det här är England , finns biljard , spelkort , schack , och badminton i balsalen . 
Avkoppling är det som står på schemat här . 
Michael , visa herrarna till deras rum , tack . 
Självklart , ma ' am . 
Den här vägen , mina herrar . 
Francy ? 
Hur länge måste jag vara här ? 
Det bestämmer tyvärr inte jag , Robert . Det bestämde er befälhavare när han skickade hit er . 
Men det kan du diskutera med dr Huston . 
Vi har bad och varmt vatten här . 
Använd det medan du kan , är mitt råd . 
Varifrån kommer du ? 
381:a . Vi flyger ihop . Och du ? 
100:e . 
När vi får chansen , kan du springa trots ditt onda ben ? 
Jag tror inte det . 
Gjorde våra pojkar det här , tror du ? 
Det verkar nyss ha hänt . RAF . 
Oj . Britterna träffade faktiskt nånting för en gångs skull . 
Okej , okej . 
Vad pågår här ? Vad gör de här ? 
Amerikaner . 
Terrorflygare ! 
Förbannade amerikaner ! 
Era jävlar ! 
Det är okej . 
Vakter ! Backa ! 
Lugna ner er . 
Sluta ! Skydda dem inte ! Låt dem klara sig själva ! Vakter ! 
Doktor Huston ? 
Får jag komma in ? 
Jadå , kom in bara . 
- Robert Rosenthal . - Ja . 
- Hur sov ni i natt ? - Okej . 
Det kan vara en konstig omställning . 
De flesta behöver ett dygn eller två . 
Det var det jag ville prata med er om . 
Jag tror inte att den här miljön hjälper mig . 
Jag vill återvända till basen . 
Varför tror ni att ert befäl sände er hit ? Vad sa han till er ? 
Jag vill veta vad ni tror . 
Det var ett uppdrag till Münster . 
Det var tufft , men jag är okej . 
Tre uppdrag era första tre dagar . 
Hundratjugo man dödade på en eftermiddag . 
Jag var inte en av dem . Jag är okej . 
Det är tredje gången ni använder ordet " okej " . 
Ni tänker inte låta mig åka , va ? 
Jodå . Om fem dagar . 
Tack , doktorn . 
" Som är i himlen , helgat varde ditt namn ... Tillkomme ditt rike , ske din vilja på jorden såsom i himlen , ty riket är ditt och makten och ... " Jag söker efter ett ställe att begrava de hundarna . 
" Och inled oss icke i frestelse utan fräls oss ifrån ondo ... " En av dem lever än . - " Fader vår ... " - Gör slut på honom . 
Klaus . Här är ett bra ställe . 
Bra . Jag kommer . 
Hjälp mig att gräva . 
Titta , en kommer visst undan . 
Låt honom gå ! Han kommer inte långt ! 
Den enskildes frihet mot en tyranns godtyckliga auktoritet . 
Detta är vad Magna Carta , eller Det stora frihetskontraktet , lade grunden till . 
Det undertecknades 1215 och är fortfarande en viktig symbol för frihet . 
Det tog förstås 500 år till för er amerikaner innan er nations grundare satte något liknande på pränt . 
Och nu i krigstid finner vi att vårt kollektiva ... Om vi inte hade varit under er kungs tyranni i 500 år , hade vi nog fått fram det tidigare . 
Vi måste vara rigorösa i våra granskningar av tidigare konflikter och hur dessa konflikter löstes . 
" Det är trevligt med en liten brasa . 
Det blir kallt där uppe . " 
- Kapten Crosby , antar jag ? - Herregud . 
Bara lugn , jag har sett män i mycket mindre , kapten . 
Stor familj , litet hus , få dörrar . Och du är ? 
Subaltern Wesgate , din rumskamrat . 
Kära nån . 
- Du väntade dig en man , va ? - Nej , jag bara ... Det var ... 
Ja , det stämmer . Ursäkta , jag väntade mig en man . 
Vi flyglottor uppmanas att dölja våra feminina namn , därav A M Wesgate . 
A står för Alessandra ... eller Sandra och M står för mitt mellannamn som jag vägrar avslöja . 
- Vi bör anmäla problemet till ansvariga . - Det behövs inte för min del . 
Jag ser att du är gift . 
Jag hoppas att din fru lärt dig att lämna toasitsen nere . 
Jo . I spegeln , var det Tracy eller Gable ? 
Det var Tracy . 
Jag gissade på Gable . 
Upp med dig . 
En kille vände sig till mig och sa : " Sir , det finns tre problem med de jädra amerikanerna . " Ursäkta språket . Han sa : " De är översexualiserade , överbetalda , och överallt . " 
Kapten Crosby . Vad säger amerikaner är problemet med oss britter ? 
Behövs inte . Nu minns jag . 
Vi är undersexualiserade , underbetalda och under Eisenhower . 
Ni amerikaner är mer rakt på ifråga om det motsatta könet . 
Som unga män skulle vi inte drömma om att pippa en debutant . 
Vi riktar in oss på kammarjungfrur och barservitriser . 
De här amerikanerna skulle bjuda en hertiginna i säng innan han tar henne ut på middag . 
Där måste jag säga emot , med respekt . 
Kammarjungfrur och barservitriser kan inte säga nej till sina arbetsgivare , men amerikanska män är ihärdiga oavsett samhällsklass . 
Och ursäkta språket , men de skulle nog " pippa " allt som rör sig . 
Det är mer än er behandling av våra kvinnor . Ni spottar på gatorna , blir stupfulla , muckar gräl i våra pubar . 
Om ni lärde era mannar lite moralisk disciplin , skulle de inte jämt bete sig som om de är hemifrån första gången och slår runt . 
Med respekt , sir , varje dag kan vara deras sista chans att slå runt . 
Så jag tänker inte mästra dem innan de får sin helgpermis . 
Du är inte stursk nog att vara pilot , men du är kapten . Så vad är du ? Navigatör ? Bombfällare ? 
Navigatör . 
Exakt vad gör du , subaltern Wesgate ? 
Lova att inte skvallra . 
Jag lillfingerlovar . 
Jag vet inte riktigt vad det är , men det låter officiellt . 
Jag är en stakare . 
Just det . 
Vad är det ? 
Jag har stakat sen min tid i Cambridge . 
Verkligen ? 
Har du gått på Cambridge ? 
Men de ger inte examina till kvinnor , otroligt nog . 
Vad läste du ? Frånsett stakning förstås . 
Nej , bara det . Vi är specialiserade . 
Var försiktig ! 
Kära nån . 
- Hur gick det ? - Ingen fara . 
Amatörer . Det tog mig flera år att lära mig staka . 
Det sitter i handleden , grabben . 
Du har aldrig stakat förut , eller hur ? 
Vad avslöjade mig ? 
Du ljuger väldigt illa . 
Ge mig lite tid . Jag ska bli bättre . Jag lovar . 
Det är inget positivt . 
Du sover visst bra än . 
Ni sa att det tar ett par dagar att vänja sig . 
Var är er ursäkt ? 
Kan inte läkare ha mardrömmar ? Visst . 
Varför inte ? 
Ni har en del bra skivor här . 
- Får jag lägga på nån ? - Visst , varsågod . 
Jag kan inte musik . Jag bara jobbar mig genom samlingen . 
Den här ... är vad ni saknar . 
Spelar du ? 
Nej . Inte alls . 
Min mor och syster fick musiktalangen , men jag vet vad som låter bra . 
Var är ni stationerad ? Norfolk . Jag är flygkirurg vid 96:e . 
Er grupp var med oss vid Bremen-uppdraget . 
Vi miste tre bombplan . 
Var det ert första uppdrag ? 
Jag miste en god vän . 
Hans första uppdrag också . 
Det här kriget ... Mänskliga varelser borde inte bete sig så här . 
- Eller hur ? - Nej . 
Men när man ser folk bli förföljda , underkuvade , måste man göra nåt , eller hur ? 
De kan ju inte strida själva . 
Så , vad ska vi göra ? Ni har rätt . Vi måste göra nånting , och här är vi nu . 
Nej , nej . Jag menar det här . Det här är precis vad man inte ska göra . 
Krocket . Rida med hundar , vad nu det är . 
Det är rävjakt . 
Man rider inte ut på rävjakt . 
Och man pratar inte om det eller klagar över det . 
Man fortsätter och gör klart jobbet , förbanne mig . 
Jag hade funnit rytmen , ni vet ? 
Tre dagar , tre uppdrag , tre hjul nere . Pang , pang , pang . 
Som Gene Krupa . 
Man stoppar inte Gene Krupa mitt i ett trumsolo , eller hur ? 
Eller två veckor senare ber honom fortsätta precis där han var utan att tappa takten , eller hur ? 
Kanske inte . Men Gene Krupa måste tänka på mer än att hålla sin egen rytm . 
Han är ansvarig för hela bandets rytm , eller hur ? 
Har aldrig druckit det rent förut . 
I Skottland anser vi att whisky aldrig ska blandas ut . 
- Skål . Okej . - Skål . 
Stor familj . Om man inte dricker ur , gör nån annan det . 
Håller du kontakten med din familj ? 
Jag är usel på att skriva brev . 
Jag åker hem när jag kan . 
Geografiskt bor de mycket närmare än din familj . Men de känns ändå väldigt långt bort ibland . 
Ja . Det är så mycket man inte kan berätta för dem . 
Dels får vi inte , - och även om vi ... - Hur skulle de kunna förstå ? 
Bara lite . Jag är inte van vid sprit . 
Senast slutade jag på golvet i ett hotellrum utan kängor . 
Berätta . 
Tja , vi var i London på helgpermis , och Bubbles kom på ett spel med småmynt och kängor . 
Jag slutade utan varken småmynt eller kängor . 
Jag menar ... Alltså . Efter det blir historien lite suddig . 
Det sista jag minns är att jag spydde på toan med Bubbles , och det fanns bara en toastol . 
- Låter väldigt romantiskt . - Jag ska väl flytta det här . 
Är Bubbles en nattfjäril ? 
Nej , nej , han är min bästa vän . 
Bubbles är bara ett smeknamn . 
Vi behöver alla nån att spy med , skuldra vid skuldra . 
Han måste vara en god vän . Ja , det var han . 
Han sköts ner i förra veckan . 
- Jag beklagar verkligen . - Det var därför jag skickades hit . 
Få komma bort ett tag . 
Det var mitt fel . 
Hur då ? 
Jag ersatte Bubbles som bombgruppsnavigatör . 
Om han hade planerat uppdragen , hade kanske inte alla de där planen skjutits ner . 
Bubbles kanske hade levat än och ... Nej . 
Din vän var ombord på planet av ett enda skäl : Att Adolf Hitler och hans banditgäng vill styra över världen . 
Inget annat . Det är enda skälet till att nån dör i det här kriget . 
Nåja , det har varit en lång dag . 
Ska vi säga god natt , då ? 
Major Egan , kom in . 
Jag är er förhörsledare , löjtnant Haussmann . 
Varsågod och sitt . 
En whisky ? Ja tack . 
Skål för potatisskörden . 
Den känner jag inte till . Skål för potatisskörden . 
Så , var ska vi börja ? 
Kanske där jag var i en stad och nån sköt de fyra som var med mig . 
Herregud . Vilken stad då ? 
- " Rüssheim , " nånting ... - Rüsselsheim . 
Tragiskt . Jag lägger till det i rapporten . 
Era kollegor , de som dödades , om ni ger mig deras namn och rang , - så kan jag vidarebefordra ... - Jag vet inte deras namn . 
Vi råkade bara hamna ihop . 
Alltså , jag uppskattar drinken och skulle uppskatta en tjockare filt , men det enda ni får veta av mig - är namn , rang , och serie ... - Och serienummer . 
Ert är O - 399510 . 
Ja , jag vet redan det . 
Samt att ni föddes i Manitowoc , Wisconsin . 
Gift ? 
Av vad jag hört , definitivt inte . 
Skvadron , 418:e . 
Grupp , 100:e bombgruppen . Tunga bombgruppen . Stationerad i Thorpe Abbotts . 
Gillar ni baseball , major ? 
Knappast en nationell hemlighet . Cigarett ? 
De är tyvärr inte lika goda som era amerikanska märken . 
Lucky Strike är min egen favorit . 
Baseball är lite av en gåta för mig , med slagträn och baser och springa i cirkel . 
Ett stort mästerskap ägde rum i förra veckan , va ? 
Ja , World Series . Just det , World Series . 
New York Yankees mot St . Louis Cardinals . 
Ett omspel , eller hur ? 
Vi ledde med 2 - 1 i matcher när jag störtade . 
Så ni håller på Yankees ? 
Vill ni veta utgången av World Series ? 
Höll Buck Cleven på Yankees ? 
Han var visst en skicklig pilot . 
- 8 : - E FLYGFLOTTILJEN KROSSAR BREMEN Jag läste om hans bedrifter vid Regensburg - anfallet . 
Han var er vän , eller hur ? 
Vi verkar skjuta ner alla era skickliga piloter . 
Visste ni att bara ett av era plan återvände efter anfallet mot Münster ? 
Ett . 
Men tillbaka till er , major Egan . 
Jag måste tyvärr säga att ni , som ni brukar säga , sitter i smeten . 
Vi vet att ni ursprungligen greps nära Ostbevern men ni finns inte listad som besättningsmedlem i nåt av planen som anföll Münster . 
Enligt Gestapo gör det er till spion . 
Då tar de fel . 
En sak kan jag tala om , major , Gestapo tar aldrig fel . 
Så jag behöver verifiering av er grupp , er skvadron och ert plan , så jag kan bekräfta för dem att ni verkligen är den ni påstår . 
John Egan . Major . 
O - 399510 . 
Major får jag säga att ni inte gör det lätt för er ? 
Gestapo är inte som jag . 
Jag är som ni : en flygare , en hederns man . 
Och jag kan förstå saker som kanske mina kollegor i de högt indoktrinerade säkerhetsstyrkorna inte förstår . 
Jag skulle vilja prata med er om Buck Cleven , John men jag vill även att ni pratar med mig . 
Om antalet nya B - 17 som väntas till Thorpe Abbotts nästa vecka , till exempel . 
John Egan . Major . O - 399510 . 
Jag förstår . 
Kaffe ? 
Hemskt gärna . 
Men skvallra inte . 
Jag kan ju inte ge alla pojkarna frukost på sängen . 
Jag ska aldrig säga nåt . 
Roligt att du har sovit . 
Jaktplan klockan tolv . Skjut ner dem , Farsan ! Kör ! 
Öppna eld ! 
In med er ! Nu ! 
In med er ! Nu ! 
Kom igen . Sätt fart . 
Jag kan inte komma över hur allt i den här stan är så gammalt . 
Delstaten jag kommer ifrån grundades 1846 . 
Den är inte ens 100 år . 
- Vilken delstat är det ? 
- Iowa . Iowa . Nog fanns det saker där före 1846 . 
Inget som ännu står kvar . 
Ja , vi får se vad som står kvar här när kriget är över . 
Finns det ett skäl till att du vägrar tala om din tjänst och stationering ? 
Ja . Och om jag hade velat tala om jobbet ikväll , kapten , hade jag gått till sherrytimmen med professor Goodhart . 
Det verkar vara en fest . 
Ska vi undersöka ? 
Mina damer och herrar , miss Ella Walsh . 
För Bubbles ? 
För Bubbles . 
Ska du inte komma in ? 
Har du glömt att vi delar rum ? Ja . Det glömde jag visst . 
Subaltern , vi har letat överallt efter er . 
Brådskande meddelande . 
Vad står det ? 
Jag måste ge mig iväg . 
- Va , nu ? - Just det . 
Ring mig när du är i London nästa gång . 
Vi går ut och dansar . 
Om du har tur , kanske jag lär dig staka . 
Det sitter visst i handlederna . 
Dina saker , då ? 
- Dem skickar de . - Det där är inte din cykel . 
Jag lånar den . 
Nöden har ingen lag . 
Sover du aldrig ? När vi har vunnit kriget ! 
- Där har vi honom . - Hallå . 
Vad förskaffar oss den äran ? 
Vi ska snart härifrån , och jag är ute efter dina pengar . 
- Oj . - Oj , Rosie . Storspenderare . Det här är killen jag berättade om . 
Berättar han historier igen ? Ja , jag har en historia . 
Vårt sista uppdrag över Münster . Vi ser alla störta , tills vi är ensamma kvar i luften . 
Ett lätt byte . 
Vi vet att de kommer för att skjuta ner oss när som helst . 
Då hör vi det . 
Är det så jag låter ? 
Vi väntar på att bli skjutna i småbitar , när den här killen , den här galna jäkeln , börjar nynna Artie Shaw . 
Helt oväntat . Det var jättekonstigt . Men jag måste säga , när jag hörde hans röst över radion var första gången jag inte kände mig vettskrämd . 
Fast han uppenbarligen hade blivit helt jävla galen . 
Jag visste att jag inte var ensam . 
Ingen av oss var ensam . 
Kom igen . Vem ger ? 
Jag ska berätta om vårt senaste uppdrag . 
Vi linkade hemåt över Kanalen , sönderskjutna , med två motorer . 
Nån anropar flygtornet på radion : " Hallå , Lazy Fox . 
G för George anropar Lazy Fox . 
Ge oss landningsinstruktioner , tack . Piloten " ... " Och andrepiloten är döda . 
Två motorer flöjlade . 
Vi har brand i radiorummet . Vertikala stabilisatorerna trasiga . 
Inga klaffar , inga bromsar , inga fallskärmar . 
Bombfällaren flyger planet . 
Ge mig landningsinstruktioner , tack . " 
Flygtornet hör det här , slår sina huvuden ihop och tänker . De tänker så fort de kan , för planet håller sig inte i luften länge till . 
Chefen för flygkontrollen tänker och tänker , tills han kommer på svaret . 
Han anropar på radion och säger : " Jag hör er , G för George . Här är era instruktioner . 
Upprepa sakta efter mig : 
Fader vår som är i himlen , helgat varde ditt " ... - Snälla . - Ni ville ju höra den igen . Vi vill inte höra det igen , så släpp det . 
Har du hört det förut ? Massor av gånger . 
Vi drog en massa olika historier . 
En del var sanna . De flesta var det inte . 
Det spelade ingen roll . 
Rövarhistorier , musik , skratt , god irländsk whisky ... Vi behövde alla nåt som hjälpte oss klättra upp i planet igen och flyga uppdrag igen . 
Jimmy ! Klarade Frankie sig ? 
Bucky ! Här borta ! 
Crank ! 
Du klarade dig ! 
Murph ! 
Glen ! 
O ' Neill , då ? 
Hallå ! Vet nån om Buck klarade sig ? 
Vadå ? 
- Jag frågar om Buck ... - John Egan ! Klockan två . 
Varför dröjde du ? 
Välkomna till Stalag Luft III , pojkar . 
Ni skulle hellre vara hemma hos era fruar . 
I NÄSTA AVSNITT Om du och jag skulle försöka rymma ? 
Min plan är att komma hem till Marge helskinnad . 
Du kan dö här helskinnad . 
- Hallå ! Sluta ! - Är det vad du vill ? 
... medan allierade trupper är fast på stränderna . 
God morgon , mina herrar . Jag är kapten Robert Rosenthal . 
Välkomna till 100:e . 
Rosie är den bästa pilot jag sett flyga en B - 17 . 
Be till Gud att du kan flyga hälften så bra som han , så kan du också klara 25 . 
De struntar i om vi alla dör , va ? 
Bra att visa de nya killarna att man faktiskt kan klara 25 . 
