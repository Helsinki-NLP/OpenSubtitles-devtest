Testar . Ett , två . 
Ett meddelande till alla boende . 
Fram till kl. 18.00 idag genomförs vapenövningar på basen . 
Det leder till en del damm och oljud . 
Trots att det kan störa de boende är träningen viktig för landets försvarsstyrkor . Ha detta i åtanke . 
De som beträder området utan tillstånd under pågående träning kan utsätta sig för livsfara . 
Alla som befinner sig i närområdet uppmanas att evakuera till en säker plats snarast möjligt efter att ha hört denna sändning . 
Det här är det bästa fiskevädret . Eller hur ? 
En kall kopp makgeolli skulle sitta fint nu . 
Grupp 1 , Lag 1 , Lag 2 . 
Kaninjakten inleds . 
950 meter till kaninen . 
Vad fan . Varför tjatar båda sidor ? Det är distraherande . 
Jinman Jeongs patetiska familjeporträtt . 
Du har haft ditt roliga . Din lögnaktiga jävel . 
Fokusera . 
Hör på , Jian . 
Löjligt . 
Kan de inte träffa från nån sida ? 
Nej . 
Huvudkaraktären utnyttjar de döda vinklarna väldigt bra . 
Ja . Filmen är slut om huvudkaraktären dör . 
Jian Jeong . Säg mig ... Här och nu , kan du se allt perfekt ? 
Ja , självklart . 
Det är uppenbart ... 
Hör på , Jian . 
Du är ingen trollslända . 
Det mänskliga ögat ser inte allt . Missta dig inte . 
Det finns alltid döda vinklar . 
Om du utnyttjar de döda vinklarna som i filmen , kan du överleva en korseld . 
Döda vinklar . 
Jian . Vad gör du ? 
Vad i helvete ? 
Lilla flicka . 
Du har sett för många filmer . 
Synd . Jag är för långt borta . 
Vad håller du på med ? 
Fan . 
De kommer från vänster . 
Diagonalt ? 
Ljudet kom från mycket högre upp och längre bort . 
Va ? 
Vart tog hon vägen ? 
- Du , Bongo . - Ja ? Kör fram en bit . Uppfattat . 
Vad gör du ? 
Ska du hoppa därifrån ? 
Ett . 
Två . 
Helvete . 
EPISODE 1 MURTHEHELP Hallå , lägg av ! 
- Släpp mig ! - Kom igen . Ta det lugnt ! 
- Kommissarie . - Ja ? Vet du vad som hände ? 
Det var jag som fick stryk . Hon spöade mig ! 
- Va ? 
- Jag är offret här ! 
- Upp ! - Lugn ! Upp och sparka mig som innan ! 
Du är för uppjagad . Var snäll och lugna ner dig , okej ? 
Ursäkta , när får jag gå ? 
Vi ska titta på övervakningsfilmerna . 
Du får gå efter det . 
Men ... - Slog du honom ? 
- Hon slog mig ! 
- Lugn , så vi hör dig . - Vad är problemet ? Låt lagen straffa henne . 
- Lägg av . - Inte ? 
Vad är det här ? 
Får jag inte gå nu ? 
Jag gjorde inget fel . Han gick in på damtoaletten . 
Jag säger inte att du gjorde något fel . Men man kan inte bara slå folk så där . 
Du skulle ha låtit bli . Du borde ha hållit fast honom istället . 
Han vill anmäla dig för misshandel . 
Han försökte slå mig först . 
Jian , du kan inte lösa det här på egen hand . 
Ring dina föräldrar och be om hjälp . Kanske en annan familjemedlem ? 
- Hej , farbror . - Jian Jeong ? 
Vem är det ? Jinwoo Park , från Yecheong-polisen . 
Jag skulle precis ringa dig . 
Va ? 
Jo ... Bli inte för upprörd . Jinman Jeong är död . 
Varför galler på femte våningen ? 
Bara en galen tjuv skulle klättra hit för att stjäla något . 
- Jag har inga pengar . - Sådär , klart . 
Och skåpet ... 
Tack för inköpet men det är inte riktigt min smak . 
Det passar inte en 20-årig tjej . 
Det är retro . 
Ni ungdomar gillar retro . 
Otroligt . 
Titta här . 
Det är gjort av järn . 
Det är skottsäkert . Det var dyrt . 
Om det blir skottlossning . 
Det låter skottsäkert , eller hur ? 
Du är säker här inne . 
Skottlossning ? Varför ? 
Glöm det . 
Bara glöm det . 
Du , farbror . Minns du närbutiksägaren som blåste mig ? 
Han bröt armar och ben i en bilolycka häromdagen . 
Sex månader på sjukhuset . 
Jag vet inte vad olyckan gjorde med honom , men han ringde och sa att han skulle betala all lön . 
Till de deltidsanställda också . 
Galet , visst ? 
Jag var så arg då . 
Jag gjorde som du sa och ropade ditt namn tre gånger . 
- Jag tror att det funkade . - Ja . 
Jag gjorde det . 
Jag bröt hans ben . 
Farbror . Du har många ärr i ansiktet , precis som en brottsling . 
Skoja inte så där . 
Varför tar du bilder på det ? 
Du går för långt . 
När en soldat faller i krig , sätter de hans id-bricka mellan tänderna för identifiering . 
Id-numret följer en från födelse till död . 
Numret är alltså väldigt viktigt . 
Vad snackar du om ? 
Det är samma sak med ditt student-id . Glöm aldrig ditt nummer . 
2-2-0-1-9-0-7-4 . 
Har du memorerat det ? 
2-2-0-1-9-0-7-4 . 
2-2-0-1-9-0-7-4 . 
2-2-0-1-9-0-7-4 . 
Det sista han sa till mig var mitt id-nummer . 
Jag undrar ... Du är Jinmans niece , eller hur ? 
Jag är vän med Jinman . 
Vi var skolkamrater . 
Du och jag träffades när du var liten . 
Minns du mig ? 
Hejsan . Hej på dig också . 
Wow ! Du har blivit så stor ! 
Så du pluggar i Seoul . Besöker du din farbror ? 
Hur mår Jinman ? 
Han är död . 
Håll inte begravningen här . 
Det andra stället är bättre . 
Det här stället är stort , men uselt . 
Jag ringer en vän som jobbar där . 
När du har bokat rummet ... 
Här är mitt kort . 
Ring mig . 
Oroa dig inte . 
Tack . 
Vi ska nu fastställa identiteten . 
Är det här Jinman Jeong ? 
En fråga ... Vid självmord , brukar inte folk skära upp handlederna ? 
Han var ensam . Hur skar han av sig halsen så där ? 
Ja , vi utredde det som misstänkt mord med tanke på skadorna , men ingen syntes på säkerhetskamerorna vid huset på en vecka . 
Enligt obduktionsrapporten kan det vara självförvållat , att döma av vinkeln på såret . Så vi drog slutsatsen om självmord . 
Jag kan skicka dig obduktionsrapporten . 
Typiskt honom att dö så här . 
Ursäkta ? 
Hans död passar honom . 
Nej . 
Skicka inte rapporten . 
Okej , då har vi fastställt identiteten . 
Vi fortsätter med överlämnandet . 
Skriv under här , så är det klart . 
Överlämnandet är nu klart . 
... två typer av sorgdräkter . 
Traditionell och modern hanbok . 
Du kan välja mellan de två . 
Var det en ny tatuering ? 
Ursäkta ! Du får inte röka här inne . 
Förlåt . 
Jag går igenom det här igen . 
Välj sorgdräkt . 
- Här är hårnålen ... - Jag är huvudsörjande . 
Vanligtvis bär män armbanden . 
Har du några nära manliga släktingar ? 
Nej , ingen . 
Det viktigaste är den avlidnes porträtt . 
Har du en bild på den avlidne ? 
Jian Jeong ? 
Det är du . 
Minns du mig ? 
Jeongmin Bae . 
Är du okej ? 
Ja , jag minns dig . Jeongmin Bae . 
Vi kan klippa ut din farbrors ansikte så här . 
Jag pluggar IT . 
Detta är lätt . 
Jag hjälpte din farbror . 
När jag kom hem efter lumpen såg jag din farbrors annons . 
Han ville uppdatera sin webbplats för jordbruksslangar . 
Jag jobbade på den i några dagar . 
Under tiden gick din farbror bort . 
Därför var jag den sista att kontakta honom , 
och den polisen ringde först . 
Ord räcker inte ... Hur kan jag trösta dig ? 
Din farbror hittades väl i badrummet ? 
Har du städat än ? 
Nej , inte än . 
Jian . Är det för jobbigt så kan jag städa upp . 
Din farbror och jag var nära . 
Det är nog okej om jag städar . 
Jag skulle uppskatta det . 
Okej . Koncentrera dig på begravningen . 
Jag städar badrummet och går hem sen . 
Tack , Jeongmin . 
Jian . 
Jag tog med Jinmans barndomsvänner . 
Lyssna noga . Du måste gengälda det här en dag . 
Gymmet vid korsningen . 
Ägaren är ordförande för Yecheongs alumner . 
De är från Yecheongs alumniförening . 
De är från Yonghan Lee . 
KAMRAT YONGHAN Jag vet inte vem det här är . 
Du har en gäst ! 
- Kom . - Okej . Jag tar hand om det här . 
Gå och hälsa på gästerna . 
Hur mår du ? 
Jag mår bra , men ... 
Jeong . Så du dog så här . 
Vi ses i helvetet . 
Önskas något annat ? 
Vill ni ha lite pannkakor ? 
Så ni var kollegor till Jinman ? 
Okej . 
Vilket gäng oförskämda idioter . 
De borde svara på tilltal . 
Är det tvillingarna från kvarteret ? 
Jag känner alla i kvarteret . 
De är inte härifrån . 
Jinman ! 
Var Jinman skyldig honom pengar eller något ? 
Eller dejtade han Jinman ? 
Han har lipat i två dagar nu . 
Jag fattar inte heller . 
Förresten , varför tog han sitt liv ? 
Han sålde slangar på internet . 
Det gick nog dåligt . 
Han hade skulder . 
Pengar är alltid problemet . 
Så varför hjälpte du honom inte ? 
Du driver sju växthus ! 
Varför skulle jag ? 
Jag har aldrig gillat Jinman . 
För att du fick stryk av honom när du rånade yngre barn . 
- Det är inte sant ! - Jo ! 
Jinman slog ut tre av dina tänder ! Jag såg det ! 
Jinman var så populär på den tiden . 
Hallå ! Hörde ni ? 
Innan Jinman kom hem igen ledde han Mokpos Getingliga . 
Vad i helvete snackar du om ? 
Han var ingen gangster . 
Jo ! Getingligan ! 
Du vet inte vad du snackar om ! 
Det här är en hemlighet som bara få känner till . 
Ryktet säger att Jinman var en anti-Nordkorea-spion för NIS . 
Vilket skitsnack . 
Det är helt befängt . 
Han hade usla betyg ! 
Han fick bara F ! 
F , F , F , F , F ! 
NIS accepterar inte så dåliga betyg ! 
Specialanställning ! 
- Getingligan ! - Jag har rätt ! 
Era jävlar ! 
Du skräms . Vad fan ? 
- Va ? 
- Vad fan ? 
Era skitstövlar ! 
Ni borde inte prata så där ! 
Minns ni inte vad Jinman gjorde för oss ? 
Minns ni när våra pappor förlorade alla sina pengar till spelhallen i grannkvarteret ? 
Varför tar du upp det nu ? 
Din pappa blev ruinerad . 
Min pappa förlorade huset . Han kom hem och eldade briketter . 
Jag och min bror dog nästan ! 
Där och då andades jag in röken och dog nästan ! 
Där och då ! 
Jinman ? 
Det var definitivt han . 
Lämnade Jinman pengarna ? 
Jinman räddade er alla . 
Jinman , din jävel . 
Vi bodde ihop i tio år men han är en gåta . 
Rök klart så åker vi . 
Jian . 
Vi åker tillsammans . 
Hon grät inte en enda gång . 
Hon kanske inte gillade honom . 
Var de osams ? Lägg av . Hon kan höra dig . 
De är otroliga . 
Alla sörjer på olika sätt . 
Bra jobbat , Jian . 
Jag städade badrummet . 
Tack , Jeongmin . 
Ingen orsak . 
För gamla tider . 
Jag är lättad att du tar det här så bra . 
Ser det ut som att jag tar det hela med jämnmod ? 
Ja ... 
Gör du inte det ? 
Jag föraktar min farbror . 
Sättet han dog . 
Jag borde inte säga så . 
Tack . 
När jag har hämtat mig kan vi väl äta tillsammans ? 
Visst . 
Ring mig , Jian . 
Hejdå . 
Jag har redan ätit . 
Men ät du . 
Vad var så svårt ? 
Vad var så svårt ? 
Du låtsades vara så stark . 
Vad ska jag göra helt ensam ? 
Jian , jag glömde ge dig det här . 
Ska jag komma tillbaka sen ? 
Jeongmin . 
Ja ? 
Jag mår inte så bra . 
Kan du stanna en stund ? 
Tack igen , Jeongmin . 
Ingen orsak . 
Jag hade ändå inget att göra . 
Jag kan stanna längre . Okej . 
Låg den i badrummet ? 
Ja , det var nog din farbrors . 
Nej . 
Vi köpte nya telefoner när jag började plugga . 
Kan den ens ringa ? 
Det kanske var en jobbtelefon . 
Som en ospårbar telefon ? 
DU FICK 70 MILJONER WON ! VAR ÄR VARAN ? 70 miljoner ? 
Hur många slangar köpte de ? 
Jeongmin . Hur mycket ? 
Arton ... 18,7 miljarder won . 
Tjänar man så mycket på slangar ? 
Nej . 
Webbplatsen du gjorde till min farbror , visa mig den . 
Slangar för 70 miljoner won ... 
Det är över 11 kilometer . 
Som du sa , det är inte rimligt att köpa slangar för den summan . 
Men webbplatsen kanske döljer en annan webbplats . 
Det här ... 
- Den mörka webben . - Va ? 
En olaglig sida . 
Slangarna var bara en front . 
En passage till den här sidan . 
Vad är det för sida ? 
Det finns priser på vapnen här . 
Det är en sida som säljer vapen . 
Vapen ? 
Sålde han det här ? 
Min farbror ? 
Vilken galen jävel ! 
Jian , ignorera det där . 
Han är galen . 
Men ska vi för säkerhets skull , ringa polisen ? 
Jinman , det är Minhye . 
Min farbror är inte hemma . 
Kom en annan dag . 
Du måste vara hans niece . 
Jag har hört mycket om dig . 
Jag är So Minhye , Jinmans privatlärare i kinesiska . 
Är Jinman bortrest ? 
Vi har en lektion idag . 
Jag ringde , men han svarade inte . 
Som du vet informerar han alltid om ändrade planer . 
Pluggade han kinesiska ? 
Det var öppet , så jag gick in . 
Är det okej om jag väntar på honom här ? 
A SHOP FOR KILLERS JIAN 7 ÅR Jag skulle ha lagat något godare . 
Struntprat . Vi äter det som serveras . 
Kom och sätt dig . 
Ja , kom och sitt . 
Är det gott ? 
Smakar det bra ? 
Det måste det vara . Du vräkte i dig allt . 
Du är bra på det . 
- Sluta . - Det är gott . 
Så varför hälsar du inte på oftare ? 
Hur längesen var det ? 
Mamma . 
- Fem eller sex år ? 
- Sju år och åtta månader . 
Nästan åtta år . 
Herregud , lillebror . 
Du har inte besökt oss på åtta år . 
Du hörde inte ens av dig . Jag trodde att du hade dött till sjöss . 
- Fattar du ? 
- Himmel . 
Sluta nu ! 
Älskling , det räcker . 
Jinman , vill du ha mer kött ? 
Ja , tack . 
Ditt ansikte ... 
- Slagsmål ? 
- Ett litet sår bara . 
Var försiktig . Min son . 
- Du måste gifta dig . - Eller hur ! Han är en luffare ! 
Kvinnor flyr från honom ! 
- Helvete . - Sluta , älskling . 
- Jian Jeong . - Min flicka . 
Vet du vad jag heter ? 
Nej . 
Jinman Jeong . 
Kom ihåg det . 
Min älskling . 
