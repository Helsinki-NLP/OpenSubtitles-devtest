KONSTNÄRSPROFIL " Inget är mindre verkligt än realism . " 
- Är du också här , Wally ? 
- Ja , de bad mig recensera nån radiopjäs . Allan . Jag trodde du hade träning till kl 16 : 00 . 
Ja , men jag gick tidigare för att se till att du kom i tid . 
Du tar det alldeles för allvarligt . 
Det är bara min mamma . Din mamma är en begåvad konstnär . 
Hon förstår drömvärlden bättre än de flesta andra . 
Nej , tack . Min begåvade mor skulle känna lukten . 
Folk som röker känner inte röklukten från andra . 
Min mor känner lukten av allt , till och med mina tankar . 
Jag är ledsen . 
Snälla , var inte det . 
Georgia O ' Keeffe sa att inget är mindre verkligt än realism . 
Jag hoppades att vi kunde börja där . 
Vad gör en konstnär till surrealist ? 
Jag vet inte om jag skulle kalla mig själv surrealist . 
Okej . 
Vad tycker du gör en konstnär till surrealist ? 
André Breton skrev i första Surrealist Manifesto ... Men vad tycker du ? 
Jag tycker ... Jag tror det har att göra med jakten på det magnifika . 
Och vad är mindre magnifikt än att försöka definiera sig själv ? 
- Det är ... - Det jag försöker säga är att era verk försätter åskådaren i ett tillstånd ... Betty , älskar du min son ? 
För jag har aldrig sett honom så galen i någon , och jag undrar ibland vart det här är på väg . 
Det är Liz från West Third igen . Jag borde ... Jag borde nog ta det . 
Ursäkta mig . Jag kommer strax . 
- Hon vill tala med mästaren . - Tja ... Håll i dig . 
Hur går det ? 
Jag är nog för förberedd . 
Jag läste din artikel i The Brownie . " USA och vi . " Den fick mig att känna mig irrelevant och gammal . 
- Du är nog nåt på spåret . 
- Ni är inte gammal , mr Durst . 
Jag vet inte om jag kände mig gammal eller bara avundsjuk . 
Nuförtiden blandar jag ihop sånt . 
Jag önskar Allen kände så . 
Om jag vore min son , skulle jag ta dig till New York . 
Hänga i Greenwich Village . 
Sen skulle jag hjälpa dig få jobb på seriös tidning . 
Jag menar , med din talang skulle du kunna gå hela vägen , Maddie . 
- Tack . - Hal , Liz vill prata med dig . 
Fråga Louise om utställningen på West Third Gallery nästa månad . 
Då börjar hon nog prata . 
- Tack , mrs Durst . - Då så . Jag ser fram emot att läsa den . 
Jag tackar mr Durst på vägen ut . 
Mr Durst ? 
Vem var hon för dig ? 
Du ville berätta Tessies historia . Du ville berätta min . 
Du ville berätta allas historia förutom din egen . 
Tessie ? Kan du höra oss ? 
Här ... Hon är här . 
Nämen , för helvete . 
Ni ljög inte . 
- Du , Paul ? - Ja . Jag ringer in det . 
Hon är så liten . 
Om det är ett sexbrott lär det bli för mycket för mig . 
- För dig ? 
- Det är Donnelly , vi har hittat flickan ... Hur visste ni att ni skulle leta här , mrs ... Schwartz . 
Jag brukar kunna se det . 
- Att peka ut judar är en livslång vana . - Hallå ! Hon råkar ha en väldigt fin näsa . 
Vet er make att ni är här , mrs Schwartz ? 
- Jag hämtar vatten åt er . - Tack . 
Vi har bara några frågor till . 
Du borde se upp , Platt . 
... och sen försökte vi gå med i den officiella skallgången . Inget nytt under solen . Ja . De hittade Durst-flickan . 
Så snabbt ? 
Bor ni här ? - Ja . 
- Vilket nerköp . 
- Tack ska ni ha . - Vänta . 
Tills någon grips kommer ni och er vän vara nyhetsstoff . 
- Så se upp för reportrar . 
- Jag planerar inte att tala med nån . 
- Jag följer er upp . - Tack . Jag klarar mig . 
Ja . Så länge du har lera i ansiktet här i krokarna , så . 
Hejdå . Godnatt . 
Fan , Dora . Jag trodde droger fick en att tappa aptiten . 
Inte med ett sånt kök som Shell har här . 
- Okej , kliv . - Kom . Kom igen . Nån här vill bli nerbäddad med mig . 
Gå försiktigt . Jag hjälper dig . 
- Dregla inte på mig . - Okej . Jag går in . - Jag ser till att hon är okej . 
- Nej . - Jag är trött , jag vill vara ensam . - Kom nu . 
Kom . En liten puss , bara . 
- Okej . - Titta till mig senare , okej ? 
Hoppas att Shell låter dig sjunga på scenen igen . 
Jag kommer att sjunga . 
Shell låter Dora vara Dora . 
Ja , så länge Dora låter Reggie bestiga henne . 
- Så är det inte . - Inte ? Vad är det då ? 
Min röst . 
Visst , du har sjungit för honom sen du var 16 , men jag minns inga gratisdroger eller rum på Gordian förrän Reggie började gilla dig . 
- Jag kanske gillar honom också . 
Dora , det finns fler ställen där du kan sjunga . 
Eggy Woods sa att niggrer åker till Paris och sjunger . 
Kan du tänka dig ? 
- Lämna hela jäkla landet bakom sig . 
- Med vilka pengar ? Jag ska leta upp Cleopatra i min drömbok , så får du satsa på ett nummer åt oss . 
Jag spelar inte med pengar jag behöver till mina pojkar . 
Jag sitter här och drömmer om att vi båda åker till Paris tillsammans . Men du följer hellre Myrtle Summer . 
Jag har inte tid med drömmar . 
Myrtle ska hitta anständigt arbete åt mig . 
Anständigt ? 
Du vet väl att Shell betalade för hennes kampanj ? 
- Det är inte sant . 
- Visst , Myrtle Summers kämpar för folket . 
Hon bryr sig om svarta kvinnor , framförallt en svart kvinna Myrtle Summer . 
- Mamma ? - Madeline . 
Vad gör du här ? 
Milton ringde . 
Har du tappat förståndet ? 
Han har varit uppe och oroat sig hela natten . 
Ja , jag tappade förståndet . 
- Var är Seth ? - Han är på uselt humör . 
Jag måste byta om . 
Madeline , tänker du berätta vad det är som pågår ? 
Tessie Durst begravs om en halvtimme . Kan vi diskutera detta efteråt ? 
- Seth vill inte gå . 
- Vad sa du till honom ? Måste jag säga något för att han ska vara upprörd över att hans mor lämnade honom ? - Jag lämnade inte honom . - Nej , just det . Du lämnade mig . 
- Vad ... Lämnade du mig ? 
Jag förstår inte . - Milton , jag behöver pengar . Jag måste hyra nåt i några veckor för att rensa tankarna . - Pengar ? Rensa tankarna ? - Jag kan inte göra det här . 
Maddie , du ville hjälpa till att hitta Tessie Durst . 
Och du hittade henne . Mazel ! Men vad pratar du om nu ? 
Kan vi inte diskutera ... 
Vi pratar . Jag pratar , du pratar . 
- Vem är du ens när du pratar så här ? - Jag vill ta en paus så jag kan räkna ut varför jag vill härifrån . 
Men nej , det låter du mig inte göra . Du vill ringa min mor , och du vill säga till vår son att jag gjort nåt fel . 
- Jag sa inte till vår ... - Han sa inget till mig . 
Kommer du eller inte ? 
Nej . Hon dog igår . 
Jag förstår inte varför vi har begravning så snabbt . 
Så själen kan gå vidare . 
Gå vidare vart , Maddie ? 
Som många i vår stad kommer du snart märka att man bryr sig mer om de dödas själar än de levandes . 
Vet du , Madeline , du borde bära svart oftare . - Du ser yngre ut . - Mamma . Det är fascinerande att du fortfarande går framåt - men alla bakvända komplimanger du ger . 
- Sluta nu . Det var ett råd . 
Människan planerar och Gud skrattar . Jag vet vad det betyder . Du har alltid sagt så . 
Hur ska du försörja dig ? 
- Jag vet inte hur du ska ha råd . 
- Jag får väl sälja bilen . 
Herregud . 
Jag är glad att min mor inte lever så hon slapp se det här . 
- Din mor dog väl under förintelsen ? - Hallå . Jag är glad att hon inte lever och ser det upprepas i USA . 
Det är en grupp 19-åriga nazister . 
De har öppnat en filial till NSRP . 
Rabbi Korn stängde shul idag ... Milton . Det räcker . 
Maddie , jag vet att vi inte känner varandra väl . Men jag hörde att du ... du vägrade lämna min Tessie när du hittade henne , och jag bara ... jag ville bara ... 
Jag är så ledsen . Såg du hennes ... Såg du hennes ansikte , Maddie ? 
Ropade hon ... Tror du att hon ropade på sin mamma ? 
Jag var inte där . - Men du ... du var där . 
Jag får henne inte tillbaka , Maddie . Jag får henne inte tillbaka . 
Vart är du på väg ? 
- Seth . Seth ! - Min flicka ! Min flicka ! 
- Jag är så ledsen . - Varför blev min ... 
Är du här ? 
Ditt jävla as . 
Jävla as ! 
Jag har ju sagt åt dig . Jag kastar ut dig om du gör om det här igen . 
Varför är du inte i affären ? 
Jävla as ! 
Min mamma trodde , att för att få ett bra jobb var jag tvungen att se så bra ut att jag inte tycktes ha några bekymmer . 
" Alla kvinnor känner till det knepet " , sa hon . 
Du fick hela ditt liv tack vare det knepet . 
Inte sant , Maddie ? 
Kontoret för kvinnligt ledarskap ... Hon är här ! 
Vem , jag ? Vad händer ? 
Linda fick WJZ att låna oss deras utrustning idag . 
Och Patricia Murphy från The Afro ska intervjua folk från samhället . 
Intervjua angående vad ? 
Hur Myrtle har hjälpt eller inspirerat dem att eftersträva förändring . 
Det du sa under eventet igår gjorde verkligen intryck . 
Hoppas du upprepar det framför kameran idag . 
Gör det nåt om jag pratar med mrs Summer först ? 
- Jag säger till att du är här . - Okej . Jag väntar där inne . 
- Ses vi snart ? - Vi ses snart . 
Ja , jag har brevet . 
Tack . Hejdå . 
Förlåt att jag stör , mrs Summer . Jag ville bara tacka för att ni bad mig hålla tal igår . 
- Du var välgörenhetseventets stjärna . 
- Jag lärde mig av den bästa . 
Kan jag sätta mig ? 
Jag hoppades att vi kunde diskutera en heltidstjänst hos er . 
Jag har dryftat din anställning och alla älskade den idén . 
Du är ansiktet utåt till hur ett bättre Baltimore kan se ut . 
Men dessvärre uttryckte några av våra vita donatorer oro över att du skulle börja hos oss , eftersom du arbetar för mr Gordon . 
Hälften av stadens färgade arbetar för mr Gordon . 
Cleo ... Det kommer uppfattas negativt om jag anställer dig efter ditt uttalande igår . 
Som om jag köpt ditt stöd . 
Men om jag arbetar för er behöver jag inte arbeta för mr Gordon . 
Ingen lämnar en man som mr Gordon , om inte han vill bli av med dem . 
- Du gjorde det . 
- Jag arbetade aldrig för honom . 
Om du syftar på de donationer jag inte längre tar emot , så förstår du säkert varför jag behöver de här donatorerna . 
Hjälp mig bli återvald , så kommer det finnas möjligheter för dig . 
Möjligheter till vad ? 
Att göra avkall på min värdighet ? 
Vi har alla fått vänta på vår tur , Cleo . 
Jag heter Eunetta Johnson och jag är 30 år gammal . 
De flesta kallar mig Cleo , ett smeknamn för Cleopatra . 
Det är vad barnen brukade kalla mig när mrs Summer var min lärare . Hon sa att jag liknade en egyptisk drottning . 
Men idag när folk ser på mig , ser de inte en drottning . 
De ser en bartender , en bokhållare en varuhusskyltdocka . 
De ser ett välgörenhetsfall . 
När jag var liten brukade min pappa säga : " Vi drömmer inte för egen del . Vi drömmer för dem som inte är här än . " 
Och jag antar att han hade rätt , för jag har inte drömt för egen del på väldigt länge . 
Men jag har två pojkar hemma , och världen tycks ge mig ett val . Jag kan behålla min värdighet eller så kan jag försörja dem . 
Jag tycks inte kunna göra båda . 
Cleopatra , är allt som det ska ? 
Cleo , raring , om du är nervös ... Cleo ! Vad är det med dig ? Se så . Cleo , raring , vi måste ... 
Okej . Okej . En paus ? 
Cleo , jag väntar utanför dörren . 
Även om du parkerar den här , kan jag inte ta den utan er makes underskrift . 
Varför måste min make skriva under om bilen står på mig ? 
För att han är er make , mrs Schwartz . 
Två tusen femhundra . Två tusen femhundra och er makes underskrift . 
- Vad sägs om 2 000 ? 
- Tyvärr , sötnos . 
Kan du köpa den här bilen utan hans underskrift ? 
- Inte än . 
- Då måste han skriva under , damen . 
Ursäkta mig . - Har ni en telefon ? 
- Ja . Där bak . 
Tack . 
- Växeln . Vad önskas ? - Jag har blivit rånad . 
Var är ni , ma ' am ? 
Nån bröt sig in i min lägenhet . 
Jag är rädd för att gå in . Kan ni skicka hit polisen ? 
- Jag behöver er adress . 
- Ovanför restaurangen The Silver Dollar . - Var ? 
I Sandtown ? - I Sandtown , ja . 
- Jag ska försöka . Hejdå . - Tack . 
Hur är läget , Sonny ? 
- Ge mig en dollar på 325 . - Visst . 
Förlåt mig . 
- Långa Teddy . 
- Har du nåt åt gamle Charlie ? 
- Jag har Jenkins , Holmes och Brooks . - Okej . - Då så . 857 till mr Brooks . 
- Jag säger det åt honom . 
Varsågod , Teddy . 
- Var rädd om dig . 
- Tack , mr Cedrick . 
Shell Gordon är en brottsling som drivit det illegala nummerlotteriet i 20 år . 
Hans enda sysselsättning är segregation och att hålla de våra beroende av honom . 
Myrtle Summer intar en kontroversiell ståndpunkt emot det så kallade nummerlotteriet . 
Denna olagliga form av dobbel spelas huvudsakligen i fattiga svarta områden och svarta arbetsklassområden landet över . 
Mrs Summers motpart menar att lotteriet finansierar svarta småföretag , en lögn vårt rättsväsende dagligen försöker fördriva . 
De som spelar på nummerlotteriet använder det som kallas en drömbok som ett försök att översätta sina drömmar till vinnande nummer , samtidigt som de långsamt förlorar sina pengar till den lokala gangstern . 
Du , titta . Släpp in henne . 
Titta på det här . 
Jag vill visa dig . Nya modell . Ful , men dubbelt så snabb som Remsons . 
Visa henne . 
Kostar ingenting . 
Och om den går sönder ? Då skaffar jag dig en ny . 
- Allt är slit-och-släng numera . 
- Sant . Såna som Myrtle och pantrarna kan skrika dagen lång . 
Det är inte rösta eller dö . Det är banken som gäller . 
Det var det jag hoppades få diskutera med er , mr Gordon . 
Jag går , chefen . 
Jag hoppades kunna acceptera ert erbjudande . 
Komma fram från bakom bardisken och sköta era röda böcker , inte bara de gröna . 
- Vad helst ni kan tänkas behöva . - Okej . Det var goda nyheter . 
Men du håller säkert med om att en man i min ställning måste kunna lita på mitt folk . 
Ni kan lita på mig , mr Gordon . 
Mitt enda mål är att kunna ta hand om mina söner . 
- Ni kan lita på mig . 
- Då ses vi väl på Pharaoh ikväll . 
Vad gäller resten , får du bevisa det med handlingar . 
- Okej ? 
- Okej . 
Om du behöver extrapengar , ta hit Slappy för att göra ett set . 
Vi ses på Pharaoh . 
- Skepp på havet . - Jag skiter i drömnummer . En bra vadhållare säljer mer än nummer . Han säljer en dröm . 
Teddy . Berätta om skeppet på havet som jag drömt om . 
Ett tydligt tecken på ett lyckligt hushåll . 
Satsa på 395 . 
- Snacka om att ha koll ... - Mitt i prick . 
- Vad har jag sagt om att ta vad , Teddy ? 
- Mamma ! Du trodde inte att jag skulle vara här , va ? Sluta . Sluta . 
- Smyga runt som en tjuv ? - Snälla , sluta . 
- Varför ? - Snälla . - För småpengarna de ger dig ? 
- Snälla . Förlåt . Lugn , Cleo . Du har sagt ditt , okej ? - Ge honom en chans . 
- Uppenbarligen inte . Jag är trött på drömbokskiten . 
- För helvete , Cleo ! - Stå här ! 
Charlie , lämna för helvete min son ifred . 
Jag tänker inte upprepa det . 
Sätt på dig jackan . 
- Du , Teddy . Oroa dig inte . - Det här är sista gången . 
Ingen fara . Jag sköter din rutt , bror . 
Teddy , vänta ! 
Teddy , vänta ! 
Tack och lov . 
- Mrs Schwartz ? 
- Ja . Tack och lov att ni är här . 
- Konstapel Platt , konstapel Davis . 
- Tack för att ni kom så snabbt . 
Ja , ma ' am . Jag patrullerar här . Ni verkar inte höra till det här området . 
- Jag flyttade hit igår . 
- Jag menar att området är fel för er . 
- Jag kan inte se er bo här . - För att jag är judisk ? 
Nej , ma ' am , inte direkt . 
Jag blev varnad , men jag trodde inte jag skulle rånas . 
Så klart . Vad är det som saknas , mrs Schwartz ? 
Smycken , främst bijouterier . Jag hade en diamantring som är borta . 
Konstapel Davis , kan du kolla om grannarna såg nåt ? Jag följer mrs Schwartz till hennes nya lägenhet . 
Tack . 
Här . 
Jag har sett er tidigare . - Men inte här . Varifrån flyttade ni ? 
- Pikesville . 
- Pikesville . - Nu bor jag här . - Stor begravning där idag . - Ja . Det kanske var där ni såg mig . 
- Är ni damen som hittade Tessie Durst ? - Det är jag . 
Och nu har ni blivit rånad . 
Det ena har säkert inget att göra med det andra . 
Det finns inte så många manikyrställen här , va ? 
Det är ingenting , bara lite smuts från flytten . 
Jag måste ringa in rånutredarna . 
Jag har ingen telefon . 
Och jag har ingen radio . För att jag inte ... Jag saknar radio , men jag har en nyckel till telefonautomaten inne på The Silver Dollar . 
Jag ringer därifrån så kan vi vänta där nere . 
- Vi vill inte röra nåt , mrs Schwartz . 
Skall vi ? 
- Tack . - Varsågod . 
- Vad snällt . 
- Det var så lite . 
En kort sekund var ni och er vän misstänkta . 
Var vi ? 
Konstapel Bosko trodde det var ett lesbiskt sexbrott eller något . 
- Ni måste skämta . 
- Jag lovar , det gör jag inte . 
Men sen hittade de akvariegrus under hennes naglar . De kommer gripa nån snubbe i fiskaffären . 
Vissa säger att de såg Durst-flickan gå in dit . 
Stackars barn . 
Får jag ställa en fråga ? - Visst . 
- Var ringen försäkrad ? 
Ni vet att det kan dröja månader innan försäkringspengarna kommer ? 
Ha det i åtanke om ni räknar med pengarna . 
- Om jag räknar med pengarna ? 
Hursom . Rånutredaren borde vara här nu . 
Kom . 
Ursäkta . 
När jag var i Memphis , hängde jag med kungen . 
- Vilken kung ? 
- Inte Martin Luther King . Elvis . 
Och jag var inte underhållningen . Vi umgicks . Jag var hemma hos honom . Jag har sett hans bilar . 
Hans barn hoppade hage . Jag frågade : " Hur gammal är din dotter ? " Han sa : " Det är inte min dotter . Det är min fru . " Jag liksom : " Åh . " 
Är allt bra ? Han är okej . 
Skräm mig inte så där . Komma hit med den där minen . 
Du blandar ihop mina miner . Det här är min " inte sitter niggern här och dricker bort dagen - när han borde söka jobb " - min . 
- Söka jobb ? Jag jobbar nu . - Jobbar ? - Så här jobbar jag . Hur många gånger måste jag säga det ? 
- Skitsnack . 
- Lägg av . Jag observerar . Sen skämtar jag om det . 
- Jaså ? - Jag kan inte jobba och skriva samtidigt . - Det vore galet . - Visst . Fattar du ? 
- Vad händer , George ? - Läget ? 
Vad händer ? 
- Ge mig två . Tack . Det här är min fru . 
- Blås röken ... Blås den ditåt . 
- Du är så rolig . 
- Jag har ju sagt det . 
Jag har fixat dig ett set på Pharaoh . Imorgon kväll . 
Hur klarade du det ? Shell . Han vill inte se ännu en svart man misslyckas . 
Men han är okej med att styra dem ? 
- Så är det inte . - Vad måste du göra ? 
- Inget . 
- Var ärlig . 
Kom igen . 
Du kan väl bara gå förbi imorgon och köra ett nytt set för grabbarna ? 
Snälla . 
Har du bytt tvål ? 
Slap , jag försöker bättra oss . 
Du måste hänga på . 
Dig hänger jag på när som helst . Fan , nu om så är . 
Kom igen . 
Värst vad du är fin . 
- Är hon inte vacker , hörni ? - Sluta . Kom . Du ser lite spänd ut . 
Vi borde göra sånt här oftare . Du luktar gott . 
För att jag är renhårig . 
Madeline Schwartz . Jag är Bob Bauer . Från The Star . 
Jag känner till er spalt . 
- Jag gillade sketcherna av er fru . - Tack . Ursäkta ... Får jag komma in ? 
Jag behöver ett glas vatten . 
Tre trappor är tufft för en tjockis som jag . 
Jag skulle inte kalla er tjock . 
Jag vet inte vad annat man kan kalla mig . 
Jag gick nästan till den andra adressen , min källa rättade mig . 
- Er källa ? - Ja . 
- Varsågod . Nån jag känner ? 
- Det kan jag inte avslöja . 
Jag lovar att jag kommer vara lika diskret med ert namn efteråt . 
Jag har dessvärre inget att erbjuda er annat än vatten , mr Bauer , och jag är inte intresserad av publicitet , så ... 
Jo , men anser ni inte att historien om hur ni och er vän fann Tessie Durst är värd att berätta ? 
Inte alls . 
Jag var också reporter en gång . 
Min make är advokat . 
Vet er make att ni och er älskare är misstänkta ? 
Jag tror att er källa felinformerat er . 
Vi är inte älskare och vi är inte misstänkta längre . 
Vem är det då ? 
- Du vet , vi betalar för bra ledtrådar . 
Om ni verkligen vill veta , så kommer mannen som grips för Tessie Dursts mord ha nåt att göra med det akvariegrus som hittades under hennes naglar . 
Ni kanske ska fråga er källa om det . 
Ska bli . 
Förresten , tack för vattnet . 
Betyder det här det jag tror ? 
Jag hörde vad som hände på mrs Summers kontor igår . Bravo . 
Det är dags för Cleopatra att se ut som en drottning igen . 
Tack , Shell . 
Stephan Zawadzkie , byggnaden är omringad . 
Låt din mor gå . 
Släpp gisslan . 
Det här är inte det du vill . 
Kom ut nu . 
Du kommer inte komma till skada om du kommer ut nu . 
Ingen skjuter ! 
Gör det inte . 
Jag lovar , kommer du ut nu så kommer vi inte att skada dig . 
Kom ut med händerna uppsträckta . 
Gör det inte . 
Kom ut med händerna uppsträckta . 
Jag är oskadd . 
Allt är okej . 
Snälla , skjut inte . Skjut inte . TESSIE DURSTS MISSTÄNKTA MÖRDARE GRIPEN 
Snälla , skjut inte . Skjut inte . Det här är min son . Han kommer självmant . 
Jag gav honom en bra ledtråd . 
Du borde ha låtit honom undersöka det lesbiska sexbrottet . 
Min far hade fått en hjärtattack . 
På tal om hjärtattacker ... Kan du be din far att ge mig respit med hyran ? 
Bara tills försäkringspengarna för ringen kommer . 
Min pappa skulle bli arg över att du frågar mig . Ja . 
Eller så är jag för rädd för att fråga . 
Jag frågar honom om du röker med mig . 
Du , Reg . Bara artister . 
Bäst du är rolig , nigger . 
- Okej . Redo ? - Klockan är 21 : 00 . 
De behöver nog ett par drinkar till . 
Den kommentaren innebär att du inte tänker vara anständig . 
Du menar ofarlig ? " Kom igen , Slap . Säg inget som gör folk obekväma . " 
Okej , ja . Du måste förstå att folk kommer hit för att glömma sina problem . 
Får väl köpa dem blå kappor . 
Mitt herrskap , vi har en speciell gäst här ikväll , och det var länge sen han stod på vår scen . 
Jag vill att ni ger en applåd för Slappy " Dark " Johnson . 
Hej , hej . Tack , tack . Wow . Kul att vara tillbaka . 
Trevligt att se så många stiliga människor . 
Svarta människor med pengar . Niggers dricker martinis nu . 
Jag är fortfarande lite nervös . Jag är ju från Södern . 
Så här många välbeställda svarta personer samlade där nere skulle få byggnaden att brinna ner . 
Det skämtet gillade de inte i Tulsa . 
Det slog inte . 
Under min uppväxt i Georgia , såg jag niggrer hänga från träden på väg till skolan . 
Jag skojar . Vi gick inte i skolan . 
Tycker ni det är stört ? Varifrån tror ni vi fick våra nya skor ? 
Såg Ferdie dig gå ut ? 
Bra . 
Han har inget med det här att göra . 
Fast kaptenen älskar att få mr Gordons kuvert . Jaså , gör han ? 
Du vet den vita flickan som hittades död härom kvällen ? 
Jag hörde talas om det . 
De låste just in galningen som gjorde det . 
Hans mamma försökte skylla det på en broder som var i affären . 
Ung färgad man med en blåtira . 
En svart man med en blåtira . 
Du ... Du borde ligga lågt tills ögat läker . 
Uppfattat , chefen . 
Harriet Tubman var nog ett bra ligg . 
Lyssna . Hon fick niggrer att lämna sina hem och fly igenom skogen och riskera sina liv för frihet ? Bara ett bra ligg får en att ta såna risker . 
Är det din snubbe ? 
- Hur visste du det ? - Smög förbi ägarens hus ... - Din blick säger allt . 
Jag måste prata med dig . 
- Allt för en chans på Harriet . 
- Du måste gå ett ärende . 
Nu ? 
Vad är det här ? 
Bara en leverans . 
Du vet inte vem som skickade dig . Adressen ligger i . 
- Är det du eller Shell som frågar ? 
- Det är ingen förfrågan , Cleo . 
Du sa till mr Gordon att han kan lita på dig . Bevisa det . 
Min son går inte ens i skolan . Där tjänar han inga pengar . 
för han fick köpa skärpet . 
Vet ni hur svårt det är att be ens barn köpa ett skärp ? Hejdå . 
Sen lämnar jag tillbaka skärpet . Vi försöker få tillbaka pengarna . 
Hur är läget , Platt ? 
Jag har nog stannat för länge . 
- Som vanligt . - Vad har jag missat ? 
De har gripit killen som klippte Durst-flickan . 
- Jaså ? - Ja . 
Du ? Släpp av mig i Bottom , så pratar jag med mrs Schwartz . 
Hon borde få höra det från polisen . 
Ms Schwartz ? 
Ms Schwartz . 
Visst , informera henne , Platt . 
Vem där ? 
Jag söker Duke . 
Är du Duke ? 
Ser han ut som en sån ? Duke ! 
Vilken fin blå kappa du har . Tack . 
Sluta skrika innan du skrämmer mina fåglar , nigger . Du och de där fåglarna . Herregud . 
Det är okej . Det är okej . 
Det var inte dig jag väntade mig . 
Jag ska bara leverera det här , sen går jag . 
Bra betalt för att ringa på och hämta cash och diamanter . 
Pengar du inte får om du inte håller käft . 
Du ... Hör på ... Behöver du en drink ? - Nej . - Säkert ? 
- Men tack . - Då så . 
Hej , baby . Hej , tjejen . 
Carol . 
Titta vem som är här . 
Jag måste tillbaka till jobbet . Ursäkta . 
Lugn nu . 
Tillbaka till jobbet för vem ? 
Fortsätter du blockera dörren får du snart veta det . 
Jaså ? 
Hon är rivig . Det gillar jag . 
Du kör . 
Nej , jag är inte här för det . Jag gör bara en leverans . Nej , nej , nej . 
Du kan inte låta en kvinna köra din - 62 Corvette . 
- Jag kör . - Sätt dig ner , fyllo . 
Fan ta din bil . Vad gäller ? 
- Vad händer ? - Hallå . 
Okej , okej . Subba , du betyder inte ett skit för mig . 
Katten är borta , så råttorna dansar på bordet . 
Jösses . Har du skrivit allihop ? 
Det är bara dagböcker . 
Vissa dagböcker är litterära mästerverk . 
- Äsch . - Hört talas om Anaïs Nin ? 
Jag har läst hennes dagböcker varje kväll . 
- Hon bodde säkert inte i Pikesville . 
- Hon bor i Paris . 
Hennes dagböcker handlar om hennes privata tankar och kärleksaffärer . 
Kärleksaffärer i Paris . 
Som att köpa bagels i Pikesville . 
Jag tänker på henne konstant . Jag har memorerat lite av hennes verk . 
Jaså ? 
" Vardagligt liv intresserar mig inte . 
Jag söker endast höjdpunkterna . 
Jag är överens med surrealisterna om att man ska söka det magnifika . 
Som författare vill jag påminna andra om att såna stunder existerar . 
Jag vill bevisa att det finns oändligt utrymme , oändliga betydelser oändliga dimensioner . 
Men jag befinner mig inte alltid i det nådatillståndet . 
Vissa dagar fylls av upplysning och feber . " 
" Vissa dagar tystnar musiken i mitt huvud . 
Då stoppar jag strumpor , beskär träd , lägger in frukt , polerar möbler . 
Men medan jag gör detta känns det som om jag inte lever . " 
Vem där ? 
Konstapel Platt . 
Ett ögonblick . 
Kommer . Ett ögonblick . 
Mina föräldrar väntar på mig . 
Glöm inte att fråga din far om hyran . 
Är allt som det ska ? 
Jag var på väg att patrullera när jag såg att det var tänt . 
Så jag tänkte informera er om att de gripit den misstänkte Durstmördaren och att vi saknar ledtrådar gällande er ring . Det bådar gott för försäkringen . 
Äntligen lite goda nyheter . 
Vore det otillåtet att erbjuda konstapeln en öl ? 
Jag tiger om ni gör det . 
Sväng här . 
Det här är Myrtle Summers hem . Det stämmer . 
Snälla , gör det inte . Ni måste inte göra det här . - Snälla . - Jag tänker inte göra ett skit . 
Jag sitter här i bilen med dig och snabba Carol . 
Vi ska titta på fyrverkerierna . 
Jag försöker tjäna ihop till julklapparna . 
Skjuter du henne kommer jultomten två gånger . 
Eller hur , raring ? 
- Det är inte min grej , mannen . - Vilken nigger . Gäller det annat än diamanter och juveler drar jag mig ur . 
Sluta spotta på min fågel . 
Fan ta dig och din jävla fågel . 
Vad fan sa du ? 
Håll dig bakom den jäveln . 
Skjut honom om han inte skjuter . 
Ge mig min jävla fågel . 
Försvinn . 
Stäng dörren , nigger . Har du en stör i röven ? 
Snälla , gör det inte . Snälla . 
Håll käften , för fan ! 
