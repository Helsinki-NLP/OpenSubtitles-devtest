Brukade mr Sabich ... Det är den andra rättegångsdagen , och i rättssalen råder spänd förväntan . 
Åklagarsidans starka öppning utlovar en fängslande rättegång . 
Din jävla skitstövel ! 
Doktor , kan du beskriva vad vi ser här ? 
Skadorna efter trubbigt våld som orsakade offrets död , Carolyn Polhemus . 
Slagen tre gånger med ett smalt , tungt föremål , vilket orsakade skallskada , svår hjärnskakning , skallfraktur och hjärnbråck . 
Tryck på kraniet gjorde att delar av hjärnan rubbades för att lätta trycket . 
Är det hennes hjärna som sipprar genom frakturen ? Det stämmer . Vad som inte syns på fotona är att den också trängde genom stora nackhålet . Det är där ryggraden går in i skallbasen . 
- Var detta dödsorsaken ? - Det hade varit det , men hon förblödde innan hjärnbråcket dödade henne . 
När avled hon ? 
Enligt kroppstemperatur och grad av likstelhet dog hon mellan kl 22 : 00 och midnatt . 
Och märkena i ansiktet ? De tyder på ett fall . Hon slogs en gång i bakhuvudet , föll handlöst framåt , bröt näsan , därav märkena under ögonen och på kinderna . 
Därefter mottog hon två slag till i bakhuvudet . 
Blåmärkena i ansiktet uppstod medan hon levde . 
De dödliga slagen kom senare . 
Fanns tecken på att hon försökte försvara sig ? 
Det fanns inga tydliga försvarssår . 
Det fanns spår av svarandens hud under en av offrets naglar . 
Är det möjligt att hon klöste honom i ett försök att försvara sig ? 
Det är möjligt . Troligare är att hon var oförberedd . 
Du sa att slaget inte dödade henne , - utan hon låg där och förblödde ? - Det stämmer . 
- Hon led . - Han leder vittnet . 
- Led hon ? 
- Det kan jag inte avgöra . 
Slagen mot bakhuvudet orsakade troligen medvetslöshet . 
Kan du utesluta att hon var vid medvetande och att hon led ? Det kan jag inte utesluta , nej . 
Doktor , har du fler resultat angående ms Polhemus ? 
Ja . Hon var gravid i sjätte veckan när hon dödades . 
Fru ordförande , jag vill härmed framlägga DNA-analysen , som överenskommet mellan parterna , vilken bekräftar svarandens faderskap . 
Noterat . 
Så svaranden gjorde offret gravid ? Ja , det gjorde han . 
Det var allt . 
Mr Horgan . 
Försvarssidan ifrågasätter inte vittnet , fru ordförande . 
- Dr Kumagai ... - Ursäkta , jag är gammal och jag måste se till att jag inte har missat nåt . Du sa " ett smalt , tungt föremål " . Som jag förstår det har du inga rön om vem som svingade detta smala , tunga föremål . 
- Det finns inget att ta på . - Det stämmer . Du har inga medicinska bevis angående vem som dödade Carolyn Polhemus . 
Jag kan bara säga med absolut säkerhet att det var ett mord . 
Och inget smalt , tungt föremål eller annat mordvapen har hittats ? 
Det stämmer . 
Tack . 
Mr Molto . Fler frågor ? 
Låt bli . 
- Vi fick det vi behövde . Gå ... - Doktor , efter obduktionen , hade du tillfälle att träffa svaranden ? Ja , han kom till kontoret och krävde aggressivt att få se kroppen . 
Är det vanligt att en distriktsåklagare dyker upp så där ? 
Det har hänt , men det är absolut inte vanligt . 
Brukade mr Sabich dyka upp för att se offer ? - Nej . - Dök mr Sabich nånsin upp - för att se ett offer personligen ? - Aldrig . 
Men han kom den dagen . Hur betedde han sig ? 
- Han var upprörd , nyckfull , rädd . - Rädd ? 
Jag förstod det inte då . Men nu gör du det ? 
Jag kände att han inte bara ville veta mina rön , utan var rädd för dem . 
Det var nåt hos honom som inte stämde . 
Det var allt . 
Doktor , har du nån psykologisk bakgrund för att ställa diagnos på uppförande när det gäller upprördhet , rädsla eller nåt " som inte stämmer " ? Jag har ett förflutet med svaranden vilket gör att jag kan uttala mig om hans beteende , och hans uppförande var ovanligt . Ni har ett förflutet . Är ni vänner ? Kollegor , inte vänner . Inte vänner . Faktum är att du anser min klient vara en skitstövel . 
- Protest . - Syftar till att påvisa fördom . 
Protesten avslås . 
Känslorna blir upprörda ibland , och jag ångrar att jag sa så . 
Du har inga fördomar mot , till exempel , distriktsåklagare ? 
Självklart inte . Det är absurt . - Har du kallat mig skitstövel ? 
- Protest . 
Fru domare , om fördomar spelar in här ... Väg orden väl . 
Doktor . 
Du och jag har också grälat några gånger . 
Så blir det ibland i vårt yrke . 
Det är en väldigt grälsjuk process under hård press , och ibland lättar vi på trycket lite grann . Men jag har absolut inga fördomar mot åklagare , och jag tar illa vid mig av antydningen . 
Har du nånsin kallat Tommy Molto skitstövel ? - Protest . - Inte oftare än du . Dr Kumagai . Kanske därför du förlorade valet . - Doktor . - Försök jobba med annat . 
Just nej . Du fick sparken , - eller hur ? - Dr Kumagai . Vi måste gå . Blicka nedåt . 
Uppfattat . Han är i bilen . 
Vi hade vad vi behövde , men du kunde inte nöja dig . 
Jag sa ju åt dig att bara få Kumagai i vittnesbåset och låta honom klargöra när hon dog och dödsorsak och vem fadern till bebisen var . Men du måste pressa på . Nu har vi en rättsläkare som framstår som en kränkt - typ som bär på agg . - Vittnesmålet var viktigt . 
Den Rusty Sabich som alla känner och älskar kunde inte ha gjort det , så vi måste visa var och när han slutade vara den Rusty Sabich . 
Jag kallar det en jävla förlust . 
Det är ett fall som kommer att bygga på indicier som tillsammans blir tillräckliga bevis . Kumagai är bara den första biten . 
Rusty Sabich var upprörd , den andra biten . 
Huden under Carolyns nagel stod inte med i den första rapporten . 
Rättsteknikerna ligger efter . Kumagai tog lite längre tid på sig med den analysen . 
Rättspatologen blir nog svårare . Jeremy Buck . 
Han är nog den bäste . Jag anlitade alltid honom . Du också . 
Han är lika precis som grafisk , så det är nog bäst att ingen av er faktiskt ser på fotona . 
Bara sakligt , neutralt , utan känslor . Okej ? 
Kan vi prata lite om kroppsspråk ? 
Vad menar du ? 
Tja , det vi såg idag var inget vidare . 
Ni måste se ut som ett par . 
Juryn kommer att ta intryck av ditt kroppsspråk , och de måste se " jag älskar honom och tror på honom " , hela tiden . 
Och om massmedia tränger på som de gjorde idag , kunde du , Rusty , kanske lägga armen om Barbara och skydda henne . 
Så juryn ska tro att han är min beskyddare . 
Ja , på sätt och vis . I den situationen . 
Raymond , jag påstår mig inte kunna ditt jobb , men att förolämpa juryns intelligens är nog inte den bästa taktiken . 
Vad de kommer att läsa i mitt ansikte är troligen chock . 
Min man står anklagad för ett hemskt mord . Hur fan ska jag kunna se annat än chockad ut ? 
Rättegångar handlar ofta om att berätta historier . 
Bästa versionen vinner . 
Du är en del av vår historia , och din vrede ger oss inget lyckligt slut . 
Det är väldigt svårt för mig att vara i rättssalen och tvingas se och höra allt som kommer att sägas , alla foton som kommer att visas . 
Att jag alls är där signalerar till juryn att jag tror på min mans oskuld . 
Jag måste vara trovärdig . Men för att vara trovärdig måste jag vara sann . 
Och det kommer jag att vara där i rättssalen . 
Jag ska låta dem se min sanning . Att jag är förfärad , att jag är äcklad , och känner avsky för denna sjuka handling , att jag är kränkt av blotta tanken att mina barns far skulle kunna begå en sån handling . 
Detta är mitt livs mörkaste stund . 
Jag tänker inte låtsas nåt annat . 
Inte inför er två . Eller för juryn . 
Vi fann hudceller under naglarna på hennes högra hand , som matchade svarandens DNA . 
Vi fann även spår av saliv i offrets ansikte och på kragen till blusen hon bar . 
DNA matchade svaranden . Märkligt nog fann vi inget DNA alls på repet som hon bundits med . 
Varför säger du " märkligt nog " ? Det var noggrant gjort . Förövaren var noga med att inte lämna några bevis . Det är ovanligt med en mordplats som är så blodig och rörig och ändå så steril när det gäller bevismaterial . 
Vad säger det dig ? 
Att stor möda har lagts på att städa upp och rensa bort spår . 
Som rättspatolog med nära 20 års erfarenhet , vad hände enligt din åsikt ? 
Enligt min åsikt skedde mordet i ett anfall av raseri oplanerat följt av ett mycket noggrann , metodisk handling att binda henne när hon var död . 
Det var allt . Tack . Har du nånsin sett en kropp bunden på samma sätt ? 
Jag hade ett mordfall för många år sen där kroppen hade bundits på ett sätt som var kusligt likt detta , ja . 
Vem var åklagaren som drev mordåtalet den gången ? 
De var två , Carolyn Polhemus och Rusty Sabich . 
Förövaren i det mordfallet heter Liam Reynolds . 
- Han fälldes . - Det stämmer . De som säkrade hans fängelsedom - var Carolyn Polhemus och Rusty Sabich . - Det stämmer . 
Efter att Carolyn Polhemus och Rusty Sabich fick honom fälld hotade han att hämnas på dem . - Är du medveten om det ? 
Jag är ingen expert på konsten att hämnas , men jag antar - att döda en och sätta dit den andra ... - Protest . 
- ... skulle vara väldigt ... - Protesten godkänd . 
Vi pratade om detta . 
Åklagarämbetet har inte utrett mr Reynolds ... De har inte utrett mig heller . Det åligger inte dem att utreda nån . - De behöver inte visa på alternativ . - Han uttalade hotelser - mot Carolyn och Rusty . - Ja , det gjorde han ... 
- Det är viktigt att juryn vet . - ... ett tomt hot ... - Varför förs inte ... - ... som du inte får utnyttja . ... detta till handlingarna ? 
Ge mig nåt påtagligt , så får du tala om det . 
I annat fall , inga fler dumheter . Fortsätt nu . 
Mr Buck , du är medveten om att min klient och den avlidna - hade en romantisk relation . - Ja . När du säger att " hud hittades under hennes naglar " , menar du verklig hud , hudflagor , som om han hade blivit klöst ? 
Nej , inga synliga hudflagor . Celler . 
Om jag kliar mig i ansiktet så här , kan man finna hudceller under mina naglar ? Det är möjligt . 
Så om Rusty Sabich kysste Carolyn Polhemus och samtidigt råkade Carolyn dra sina naglar över hans nacke eller rygg , kan det inte förklara salivspåren som fanns på henne och det DNA som fanns under hennes naglar ? 
Jag antar det . Så det DNA som du menar visar att han dödade henne kunde lika gärna visa på att han kysste henne ? 
Du förstår skillnaden ? 
Visste du att svaranden och ms Polhemus hade en relation ? 
- Jag blev medveten om det . - Hur då ? 
Tja , jag hade olika skäl att misstänka det . 
Beträffande när jag visste säkert ... Jag skulle lämna av en fil på Rustys kontor . 
Det var sent . Jag trodde han var borta . Det var han inte . Jag klev in . Han kysste Carolyn . 
- Här är Roberts fall . - Ja . - Jaha . - Ja . 
- Tack . Ja . - Såja . Vi ses imorgon . Jag skyndade iväg , och hon följde efter mig . Det var otroligt pinsamt , och jag gick . 
- När var detta ? 
- I februari . 
Var du vittne till fler tillfällen ? 
Inget direkt sexuellt , bara kontorsskvaller . 
Men visst fanns det underströmmar . 
Som till exempel ? 
En gång såg jag dem i parkeringsgaraget . 
De ... Jag vet inte ... Jag tror att de grälade . 
- ... tillsammans . Jag vet inte . - Håll dig borta . Jag ställer ju bara en fråga . Kan du inte bara ... 
Men för i helvete . Hon satt i sin bil , han bankade på bilfönstret , och hon körde iväg . 
Hade du tillfälle att diskutera detta med mr Sabich ? Ja . 
Vad sa du ? 
Jag sa att jag var orolig att han höll på att , jag vet inte , gå överstyr . 
- Gå överstyr ? - För hennes skull . 
Han började gå upp i limningen , blev fixerad . 
Tyckte du inte om den här relationen mellan mr Sabich och ms Polhemus ? - Du ogillade den ? - Det stämmer . Och du ogillade Carolyn Polhemus , eller hur ? 
Det var inte det . Det var oprofessionellt . 
Du gillade inte Carolyn , eller hur ? Nej , det gjorde jag inte . 
Rapporterade du saken till personalavdelningen ? 
Nej , det gjorde jag inte . 
Och såvitt du vet gjorde ms Polhemus ingen anmälan till personalavdelningen om mr Sabich ? 
Det stämmer . 
Vet du om hon nånsin anmälde nån till personalavdelningen ? 
Ja . Vem då ? 
Tommy Molto . 
Har du kännedom om att jag skulle ha uppträtt oprofessionellt eller olämpligt gentemot ms Polhemus ? 
Jag har ingen sån kännedom , nej . 
Och har du nån kännedom om klagomålet som lämnades in ? 
Jag vet bara att hon inte ville jobba på några fall med dig . 
Hon kände sig äcklad av dig , sa hon . 
Okej . Såg du mig nånsin uppträda oprofessionellt mot offret ? 
Inte direkt . 
Rusty Sabich , då ? 
Svaranden verkade fixerad och gick överstyr för hennes skull . 
Är det ditt vittnesmål ? Det stämmer . 
Tack så mycket . 
Jag tycker nästan synd om Tommy . 
Det gjorde nästan jag med , tills jag mindes att han är en förbannad kackerlacka . 
Man kan inte mosa honom . Han kommer tillbaka hela tiden . 
Och han fick fram det han ville . 
Du är orolig . 
Tja , om juryn håller fast vid bevisbördan är jag nöjd med vårt läge , men om de behöver nån att lägga skulden på , är det Rusty . 
Allt väl ? Jadå . Och du ? 
I psykologin i skolan har vi läst om trauma och dissociation . 
Hur hjärnan kan skydda en från en själv . Som ett slags ofrivillig bortkoppling från verkligheten . 
Har du nånsin känt så ? 
Hur menar du ? 
Bara ... Folk kan fjärma sig från sina minnen . 
Om ... Om man gör nåt man inte kan förlika sig med eller hur man ser på sig själv kan det orsaka dissociation . 
Mitt minne fungerar bra . 
Rusty , jag måste prata med dig . 
Alltså , för några månader sen ungefär när jag blev avskedad från galleriet , började jag gå till en bar på dagarna . 
Och där fanns en bartender som var fil dr i konst . Vi började prata och det klickade verkligen mellan oss och vi kysstes . Jag kysste honom . 
Men det var allt som hände . 
Det var bara en distraktion . Det var ... Det var bara en kyss . 
Var hände det ? 
I hans lägenhet . 
- Jag ville se hans konst . - I hans lägenhet ? 
- Det var allt . - Du ville se ... - ... en bit av hans konst ? - Låt bli , Rusty . 
- Låg du med honom ? - Nej . 
Varför berättar du det här nu ? 
Jag vill vara uppriktig mot dig . 
Jag trodde att vi skulle vara det mot varandra . 
Jag står inför rätta ... och riskerar livstids fängelse . 
Uppriktiga ? 
Jag vet . 
Du grillar mig varenda dag . 
Du grillar mig . " Vad hände här ? " " Vad hände där ? " " Varför berättade du inte om er ? " Fråga efter fråga . 
Och när jag säger : " Jag försöker bara vara uppriktig , jag försöker bara säga vad som hände såvitt jag minns det . Jag kan inte förklara hur jag tänkte " , grillar du mig om och om igen . - Så orättvis du är . - Och igen . Orättvis ? Inte rättvist , Barbara ? Vad är rättvist ? Vad är rättvist nu ? 
Hur känns det ? Va ? 
Hur känns det ? Att begå ett jävla misstag ? 
För i helvete . 
- Dra åt helvete , Rusty . - Jag dra åt helvete ? 
- Jag går nu . - Är mina bilnycklar i köket ? 
Skölj av era skålar , tack . - Jadå . - Här är de . 
- Glöm inte geometriläxan . - Den är i väskan . - Följer du med ? 
- Nej , jag ska träffa Lorraine . - Jag är sen . - Barbara ? 
Kyle , har du din lunch ? Jadå . 
Jag kan följa med och fylla en plats . 
Raring . Det behövs inte . Det är säkert . 
Förlåt om jag gjorde dig upprörd igår kväll . 
Varför berättade du för honom ? 
- Jag vet inte , Lorraine . - Det var en usel idé . Jag vet . 
Det är bara det att vi nyligen har ... Jag tänkte ... Jag kände att vi fick kontakt igen . 
- Jag kände mig ... - Mm . ... nära honom och trygg . - Och ... - Okej . ... det där med Clifton kändes så betungande och jag behövde ... 
Ja . Och det blev inte bra ? 
Och därför ska du inte gå till rätten ensam mer . 
Jag kommer att vara med dig . 
Jag ska gå dit igen , men inte idag . 
Idag är det allt de tagit från hans och hennes datorer . Ja . Jag kan nog inte sitta där och lyssna på alla hans kärleksbetygelser ... - Herregud . - ... och så vidare . 
Vet du , kvällen hon mördades sms:ade han henne 30 gånger . 
Det är nog faktiskt det mest graverande i hela fallet . 
Trettio gånger ? 
Och pappan har just lagt in om en domstolsorder som hindrar att hans son behöver vittna . 
- Är det sant ? - Jag avslår begäran . Men jag förstår hans motiv . Den här dagen blir otroligt jobbig känslomässigt för en grabb som redan är i obalans . 
- Han är ett nyckelvittne . Så ... - Låt mig fortsätta . 
Jag vill bespara familjen mer onödig smärta , vare sig den är onödig eller inte . 
Det här fallet är som mest dråp , och det vet ni . 
Även ert eget vittne sa att det troligen var oplanerat . 
Glöm överlagt mord . Och mina instruktioner blir ingen draghjälp . 
Att du är fri mot borgen är också lite magstarkt . 
Dråp tycks som en bra medelväg . - Glöm det . - Nej . 
Ni får er fällande dom . Du får återuppta ditt liv om åtta år . 
- Det är rena gåvan . - Jag accepterar ingen dom . Nedlagt åtal och en ursäkt är det enda jag accepterar . 
Sista chansen att anta erbjudandet . 
Nån som vill backa ? 
Okej . 
Båda sidor tar det försiktigt med pojken . 
Hej , vännen . 
Vill du gå upp och lägga dig ? 
Spring upp och lägg dig . 
Minns du när de var ... När de var små och sov , satt vi och såg på dem i timtals . 
Som skyddsänglar . 
Varför stannar du ? 
Av samma skäl ... som du . 
Michael , du och jag träffades förut , så jag beklagade sorgen . Jag vill göra det ännu en gång . Både för förlusten av din mor , men också för traumat att behöva vara här idag . Det vi ber dig om är hemskt , men det är för att en mycket hemsk sak hände din mamma . Mr Molto . 
Jag vill rikta din uppmärksamhet till kvällen då din mor mördades . Kan du berätta var du befann dig ? 
Jag åt middag hemma . Jag såg på tv eller nåt . Kanske spelade tv-spel . 
Jag lämnade huset senare och åkte dit . 
För att klargöra , du lämnade huset där du bor med din far , Dalton Caldwell , och sen åkte du dit , säger du . Var är " dit " ? Där mamma bor . 
För att göra vad ? Min mamma och jag gick inte ihop . 
Hon ville inte ha mig där . 
Jag var inte välkommen . Det gjorde mig förvirrad . Ibland åkte jag bara dit för att titta . 
Titta ? 
Se det liv hon inte ville att jag skulle vara en del av . 
Jag förklarade visst det här förut . 
Åkte du till din mammas hus ofta ? Då och då . Jag vet inte . Kanske en eller två gånger i månaden . 
Vad gjorde du när du kom dit ? 
Oftast stirrade jag bara på huset på avstånd i mörkret , så att hon inte skulle se mig . 
Ibland såg jag folk gå in . Oftast han . 
Notera att vittnet syftar på svaranden , Rusty Sabich . 
Jag visste vad de gjorde . - Protest . - Bifalles . 
Svara bara på frågorna , Michael . 
Och om du känner att du behöver en paus , säg bara till , okej ? 
- Jadå . - Då fortsätter vi . Okej . 
Tog du de här filmerna ? Ja . 
Den 16 juni . 
Kan du läsa datumangivelsen längst upp i bild ? 
Ja . " Kl 21 : 49 . " 
Och återigen , var detta det du filmade kl 21 : 49 , - kvällen din mor mördades ? - Ja . 
Efter din mors död , sms:ade du svaranden ? Ja . Vad skrev du till honom ? 
Jag skrev : " Du var där . Jag såg dig . " 
" Jag såg dig " , vadå ? Vid huset när jag filmade . 
Bad du att få träffa svaranden ? 
- Ja . - Varför gjorde du det ? 
Jag ville se den som mördade min mamma i ögonen . 
- Protest . - Bifalles . 
När du hade begärt ett möte , träffades du och svaranden ? 
- Ja . - Vad pratade ni om ? 
Han frågade varför jag ville träffas , och jag sa att jag ville se den man i ögonen som mördade min mor . 
Protest . Bifalles . Vittnet uttrycker bara sin åsikt . 
Anklagade du svaranden för mordet på din mor ? - Ja . - Hur svarade han ? 
Han förnekade det . Men jag såg att han ljög . 
- Protest . - Bifalles . 
Michael , du får uttrycka dina intryck , men fastslå dem inte som fakta . Okej ? 
Okej . Pratade du nånsin med din mor om svaranden ? 
Som sagt hade vi inte mycket kontakt . 
Hon berättade inte mycket . Men cirka två veckor innan hon dog berättade hon att hon hade problem med en man på jobbet . 
Det var mitt intryck att det var samma man som hon hade en affär med . 
Sa hon nåt mer ? 
Att hon började bli rädd för honom . 
Har du nån aning om vem hon menade ? 
- Protest . Spekulation . - Protesten avslås . 
Mitt intryck var att det var samma man - som jag fick intrycket mördade henne . - Protest . 
Samma man jag tog foton av kvällen hon mördades . 
- Protest . - Bifalles . Svara bara på frågorna , Michael . Spekulera inte . 
Tack , Michael . Inga fler frågor . 
Du får många intryck , eller hur ? 
Du fick intrycket att din mamma var rädd . Du fick intrycket att det var mannen hon hade en affär med som hon var rädd för . Intryck . Det är ett märkligt ord . 
Låt oss prata om det ordet lite grann . 
Vad betyder ordet ? Det betyder tron eller övertygelsen om nåt man inte har sett , eller hur ? 
Advokaten ? 
Mr Horgan , har du en fråga ? 
- Ray ? Ray ? - Jag är hans fru . 
- Ingen puls än . - Igen . Redo ? - Tre , två , ett , undan . - Det ordnar sig . 
