Inga allierade . 
Ingen hjälp . 
Du är helt ensam , Keyleth . 
Men du har tur . 
För du får se min nya ståtliga kropp . 
Det perfekta vapnet att förstöra alla asharibyar med , en efter en . 
Det ska du inte . 
En sån formel hade kanske förstört min gamla form . Men jag har blivit döden , barn ! 
Keyleth ! 
Thordak ! 
Jag tror att det är Raishan . 
Har hon bytt kropp ? 
Jag måste inte förstå det för att döda den . 
Den här kroppen känner ingen smärta . 
Hand ! 
Kom . Med mig . 
- Pike . 
- Ska bli . Gå ! 
Nu är det slutlekt ! 
Kan inte ... Se upp ! 
Kom igen . 
Jag klarar av eld . 
De här lågorna bränner på annat sätt . 
Pikey ! 
Tror ni att jag hade hjälpt er att få tag i relikerna om de var ett hot mot mig ? 
Ni är marionetter ! 
Jag drog i era trådar och ni dansade . 
Keyleth ... Keyleth ! 
Keyleth ! 
Fly . Ge dig av därifrån . 
Jag har en plan . 
Gör inte det mot mig , Kiki . 
Gruppen tar risker hela tiden , nu är det min tur . 
Vax ... Lita på mig . 
Raishan ! Låt dem gå . 
De orsakade inte din sjukdom . 
Det var mitt folk . 
De är dina fiender ! 
Asharierna var allierade med min sort en gång . 
Tills de bedrog oss och gjorde anspråk på naturen själva . 
Du skulle göra likadant . 
Det är en lögn . 
Spela inte naiv , Keyleth . 
Du firade att ni dödade Brimscythe , Umbrasyl , Vorugal ! 
Vi båda drivs av ambition . Erkänn ! 
Bjässen , har du fler slag i handskarna ? 
Vi kollar . 
Ingenstans att fly . 
Kom igen , fortsätt . 
Farväl , barn . 
Skynda dig , Grog ! 
Nej ! 
Du tyckte om henne . 
Så synd . 
Thordak dödade din mamma . 
Då är det inte mer än rätt att han dödar dig med ! 
Va ? 
- Keyleth ? 
- Omöjligt . 
Min sjukdom ? 
Nej ! 
Du får inte ! Inte igen ! 
Du kan inte skada den här kroppen ! 
Hon verkar just ha gjort det . 
Ashari ! Snälla . Hjälp mig ! 
Jag vet inte hur du gjorde det , men du var legendarisk . 
Sjukdomar är en del av naturen . Och man kan kontrollera den om man hittar sitt ankare . 
Tänker du kyssa mig eller ? 
Vänta . 
Förlåt . Det är inte du ... Det är giftet . 
Så tjockt . 
Korpdrottningen , guida mig . 
Du har sökt mig för ett korrupt syfte . 
Är det fel att befria min vän från evig plåga ? 
Vi hedrar övergången från liv till efterlivet , vi kränker det inte . 
Hans själ är redan kränkt ! 
Om du mixtrar med döden får du känna på ännu värre sorg . 
Om du tar tillbaka honom , blir det till ett pris . 
Så det finns ett sätt . 
Visa mig . 
Visa mig ! 
Om Raishan kunde överföra sin själ till Thordak , varför kan inte vi återföra Percy till sin egen kropp ? 
Ja , men vad händer om du trotsar Korpdrottningen ? 
Hon är en gud . Okej . Något som djävulen Zerxus sa har fastnat . 
Ibland ska man gå emot sin guds önskan . 
Gudarna skapade oss inte för att följa dem blint , eller hur ? 
Vex hade varit död i några minuter när du återupplivade henne . 
Percy har varit borta ett tag . 
Han kanske blir en zombie . 
Och även om vi kan , så har hans ande lämnat det här planet . 
Nej . 
Jag har känt att hans själ hålls fången i Orthax . 
Vänta . En själ i en demon ? 
Var är demonen ? 
Okej . 
Jag behöver sprit . 
Pickle , om du återställer hans kropp , tar jag kontakt med Orthax . 
Percy dog nästan när han bröt Orthax förbannelse . Ska du göra det utan Korpens hjälp ? 
Hon varnade mig att det är farligt att utmana ödet . 
Det betyder inte att det är omöjligt . 
Vax , om du inte återvänder ... Om jag förlorar Percy och dig ... Syster ... 
Ingen kan ändra det förflutna . 
Man kan åtminstone försöka . 
Kroppen blir inte bättre än så . 
För tur . 
Orthax , jag söker hämnd . 
Mot vem ? 
Mot dig . 
Det har börjat . 
Varför har du kommit , Korpmästare ? 
Det finns inget här för dig . 
Percival De Rolo . 
Jag kräver att han släpps . 
Percy tillhör mig . 
HÄMND Det gör alla . 
Han följer inte med , även om du hittar honom . 
Släpp mig ! 
Jag kommer , Percy ! 
Det här blir mycket svårare utan Kash . 
Jag hjälper dig . 
Du kanske också hör hemma här . 
En rädd liten pojke intvingad i en pakt med Korpdrottningen . 
Du måste lyda hennes minsta vink ... Annars straffar hon dig med en hemsk framtid . 
Håll ner honom ! 
Men jag kan skydda dig från pakten . 
Du kan , precis som Percy , vara fri här , fri från hennes makt . 
Ge efter för ditt hämndbegär , mästare , för Korpdrottningens öde kan inte ändras . 
Men det kan böjas . 
Hans kropp är redo ... Men formeln håller inte länge . 
Vax . Vax ! Hör du mig ? 
Skynda dig ! 
Vad är det här för ställe ? 
Percy , guida mig . 
De Rolo , hör du mig ? 
Percy ? 
Vem är du ? 
Vi måste gå . 
Nej . 
Jag har jobb att utföra . 
Jag vet inte vad den har gjort med dig , men det här är inte du , Percy ! 
Släpp mig ! 
Jag vet inte vem du pratar om . 
Ser du ? 
En själ kan inte räddas från min domän . 
Särskilt inte en som inte vill lämna . 
För helvete ! Lyssna på mig . 
Hans skam driver min smedja . 
Eldens dån kan inte dränka hans skuld . 
Percival förtjänar det här . 
I helvete heller . 
Om du ändrar hans öde , Korpmästare , blir du aldrig densamma ! 
Aldrig att känna lycka ! 
Vakna , De Rolo ! Kom igen ! 
Vi kan inte hålla den . 
Det måste ske nu . 
- Hur ? 
- Jag vet inte ! 
Det finns ingen manual ! 
Jag vet inte om du hör mig , men dina vänner behöver dig . 
Fan , jag behöver dig ! 
Percy . 
Det var inte så här det skulle ske . 
Och du skulle avsky all uppmärksamhet , men dagen med dig i Syngorn , när du stod bredvid mig och lät mig vara del av något som du håller kärt ... 
Du stod upp för mig och jag ljög för dig . 
Och för mig själv . 
Jag var för rädd för att erkänna det . 
Du är fascinerande , obstinat och den smartaste mannen jag känner . 
Du måste hitta tillbaka till oss , Percy . 
Snälla ! Kom ihåg vem du är ! 
För sanningen är ... Jag älskar dig , älskling . 
Mitt hjärta ... Det är ditt . 
Vex ' ahlia ... Vänta . 
Tillbaka till smedjan . 
Nu ! 
Hon älskar dig . 
Och jag med ... broder . 
Nej . Nej ! 
Det är mitt rike ! 
Du tillhör mig ! 
Gör det nu ! 
Du har något där . 
Försiktigt . 
Jag har precis börjat andas . 
- Ja ! 
- Så underbart . 
Helt otroligt . 
Vax . 
Jag är här , Stubby . Jag mår bra . 
Det var en lättn ... Bättre , älskling . 
Du tog dig till porten två gånger . 
I den här takten joggar jag när jag fyller 60 . 
Så länge det där nere fungerar är det lugnt . 
Tack för allt . Särskilt för att du inte gav upp . 
Kom ihåg , jag dog också en gång . 
Jag trodde inte att upplevelsen passade en man av din rang . 
Kan ni stappla tillbaka till middagen ? 
Scanlan har kyckling på gång i slottet . 
Trinket ! Ge lorden lite hjälp . 
Vax , jag har dig att tacka för mitt liv , broder . 
Det glömmer jag inte . 
Inte hon heller . 
Han serverade åtminstone champagne . 
Du , bjässen ! Kan du skicka kniven ? 
Kompis ? 
Ja , kniv , jag gör som du befaller . 
Helvete . 
Måste döda ! 
Se på ditt dumma ansikte . 
Dummer . Du lurade mig en kort stund . 
Varje ögonblick med er är surrealistiskt . 
Du älskar det . 
Gilmore ! 
Det luktade kyckling . 
Det är vår Scanlan , han är köttmannen . 
- Hur är Whitestone , Shaun ? 
- Fantastiskt ! Lady Cassandra bjuder in er alla för att fira Vinterkrönet . 
Toppen ! 
Shopping ! 
Jäklar . Det förtjänar en skål . 
Scanlan , har du en sång för det ? 
Ja , det har jag . 
Men innan det , jag har tänkt och ... Vårt uppdrag är över . 
Och fast vi inte borde ha lyckats , så gjorde vi det . 
Men med alla skatter vi hittade och äventyret vi har haft , har jag sökt något annat . 
Jag försökte på fel sätt , men den rätta hittade mig . 
Det låter smörigt , men jag gillar mig själv bättre när jag är med Kaylie . 
Hon är betydelsefull för mig . 
Och jag tror att jag för första gången i mitt liv är betydelsefull för henne . 
Men du är betydelsefull för oss med . 
Ni är som min familj . 
Men nu har jag en riktig familj . Och hon är bäst . 
Jag vill inte dra ner stämningen . Jag ville bara säga att vi ger oss av efter middagen . 
Vart då ? 
Världsturné låter bra . 
Okej ... Det här är jobbigt . 
Jag har lagt min aramenté åt sidan . Men det är dags att bli den jag är menad att vara . 
Så vi kommer också att sticka . 
Stormens röst kan behöva en väpnare , och jag är snabb på att hämta vatten . 
Jag är glad för er skull . 
Rym inte iväg och gift er bara . 
Och oroa dig inte , Gilmore , Percy och jag följer med till Whitestone . 
Lady Vex ' ahlia har trots allt inte upplevt livet som adel än . 
Vänta lite . 
Betyder det att vi gör slut ? 
Jag försvinner inte . 
Och om fara uppstår igen , vilka tror du att de kontaktar ? 
Dråparskrået ? 
Rikets beskyddare , dummer . 
Vi är fortfarande Vox Machina . Och vi sabbar fortfarande saker . 
Ja . Det skålar jag för . 
Skål ! 
Ja ! 
Så ska det låta , bjässen . 
Jaha , pappa ? Ska vi ? 
Det är i stunder som dessa Som man ifrågasätter allt 
Typ , varför är jag här ? 
Och du där helt ensam ? 
Jag vill säga rätt saker Men jag hittar inte orden 
Jag vill bara prioritera dig DER KATZENPRINZ OCH ANDRA SAGOR 
- Jag skulle bränna mig 
- Bränna Om det betydde att jag kunde rädda dig Inte ens tveka att gå genom eld 
Om det var enda sättet att ta mig till dig 
- Jag skulle korsa världen - Jag skulle korsa världen 
- Och inte stanna förrän jag hittat dig - Hittat dig 
- Jag skulle leta efter stjärnorna - Jag skulle leta efter stjärnorna - Hoppas att de leder mig till dig 
- Jag skulle korsa världen - Jag skulle korsa världen 
Vi är hans ögon . 
Vi är hans röst . 
Vi är hans beröring . 
Vi är hans hjärta . 
Vi är hans blod . 
Vi är hans blod ! 
