Det är viktigt vad ens kläder uttrycker . 
Det är inte fel att anpassa sig , bara man vet att man gör det . 
Jag kanske klär mig som ett får , men det finns en del tecken som avslöjar för den observanta att jag snarare är en varg i fårakläder . 
- Har ni planerat när ni ska avslöja er ? 
En ny kostym för en ny era . 
Hans själ är stark , och kroppen kommer att följa själen . 
Det låter trösterikt . 
Försök hämta tröst i det . 
Jag vill inte göra nåt som förargar dig eller din far . 
Du har fria händer , John . 
Geoffrey . 
Ursäkta att jag stör , Ers nåd . Väntar ni besök ? 
Jag ser fem fordon på Field Barn Lane . 
Nej , absolut inte . 
Verkar de vara härifrån ? 
Nej , de ser inte ut som några fritidsflanörer . 
Okej . Stanna där , så kommer jag . 
" Släpp loss din vrede på de som motsätter sig ... " 
Jag kollade fågelholkar när jag fick syn på dem . 
De har varit här i 20 minuter . 
De verkar mena allvar . Vet du vem de är ute efter ? 
Det är en gudfruktig kokainlangare från Liverpool . Det här bådar inte gott . 
- Amen . - Amen . 
Freddy , har du hört nåt från Gospel-John ? 
Om jag hört nåt från Gospel ... Visst . Vi messar och utbyter tapetidéer . 
Varför skulle jag ha kontakt med den blådåren ? 
Okej . Säg åt alla att hålla sig inomhus . Visst . Men vad fan är det som pågår ? 
Jag ringer när jag vet mer . 
Vi måste hämta några saker i min stuga . 
Är det inte lite överdrivet ? 
Det är mitt jobb att döda ohyra , Ers nåd . 
Jag har gjort nåt dumt , mamma . 
Och han där ute verkar ha fått reda på det . 
Hej , Freddy . 
Jag vill driva in en skuld . Nåt som du är skyldig mig . 
Vi kan göra det här på två sätt . 
Du kommer ut , eller så kommer jag in . 
- Hej , pappa . Hur är det ? - Strunt i det . Vad är det senaste ? 
Jag har pratat med läkaren . Jack mår bättre . Han sover , men det går åt rätt håll . 
Jag pratade med Eddie och har funderat . 
Du måste komma hit på en gång . Ta med dig hertigen . 
- Det kan bli svårt . - Varför det ? Tja , han svek oss , så jag svek honom . 
Du borde ha bättre koll på nyheterna . Du verkar ligga 24 timmar efter . 
Se till att lösa det , vad du än har gjort . Jag behöver en nöjd hertig . 
Jag kan ha ringt till Gospel . 
Vad i helvete ? 
Susie , Gospel-John har precis kommit till godset . 
Förlåt för det . Det är nog mitt fel . 
Vad fan gjorde du så för ? 
Jag hade mina skäl . Är han där ? 
Han och halva brödraskapet . 
- Håll ut . Kavalleriet är på väg . - Okej , men skynda dig . 
Jimmy , lyssna noga nu . 
Hertigen är i knipa . 
Jag skickar dit några killar . Släpp in dem i huset . 
Ursäkta , John . Min bror är här . Ett ögonblick . 
Mr Dixon . Du inkräktar på privat egendom . 
Jag tänkte återlämna hagelbössan . 
- Din bror skulle få den . - Eddie , jag går ut . 
Jag ska ge er fem minuter av respekt för släktens arvegods . 
Så bra . 
Tammy och mamma , stäng fönsterluckorna . 
Nu får det vara nog . 
Jag älskar er alla . 
- Det var fint att känna er . - Freddy ! 
Nej , det är min soppa . Jag får ta smällen . 
- Du får inte . - Det är lugnt . 
Hör ni , det är lugnt . 
Jag förtjänar det faktiskt . 
Jag är en riktig skitstövel . 
Om de låter mig leva återgår jag till att vara en skitstövel . Eller hur ? 
Har jag fel ? 
Där ser du . Men det är lugnt . 
För nu kan jag för en gångs skull göra nåt osjälviskt . 
Jag kan återfå en gnutta värdighet . 
Ta inte ifrån mig det . 
Gör inte det . 
Det är inte värdighet . Det är smärta , våld och död . 
Vi älskar dig . 
Och ja , du kan vara lite av ett as ibland . 
- Ett stort as . - Ja . 
Men nu behöver vi dig . Okej ? 
Jag behöver dig . 
- Okej . - Bra . 
- Mamma , ta med personalen ner i källaren . - Ja . 
Jag hämtar Charly . 
Var försiktiga . 
Tammy , se till att dörren är låst . 
Vi tre mot en jävla gangsterfamilj ? 
Har du nån plan , Edward ? 
- Bra . Ingen plan . Först värsta talet ... - Lägg av ! Vad har du för plan ? 
- Det är helt ... - Ska du ge upp ... Ers nåd . 
Jag har fem hagelbössor till , och ett gevär . 
Perfekt . Okej . 
Det har snart gått fem minuter . Ska vi köra igång ? 
Ers nåd , vad har vi för plan ? 
- Hjälpen är på väg . - Okej . 
Det här förändrar läget en aning . 
Jimmy , vad känner du inför det här ? 
Inget för mig . Jag är pacifist . 
Okej . Källaren med mamma och de andra . 
Geoffrey , ta övervåningen . Alla andra , hitta positioner här . 
Var är mitt maskingevär ? 
Skit samma . 
Vet du varför jag älskar duvor ? 
De symboliserar harmonin mellan människan och naturen . 
Redan innan Noah gick i land samarbetade människan med fåglar . 
Har du hört talas om Cher Ami ? 
I slutet av första världskriget var 500 franska soldater fast bakom fiendelinjen . De blev beskjutna av sina egna . 
En major sände iväg en duva efter hjälp . 
Duvan blev skjuten i bröstet , förlorade ett öga och hade ett ben som knappt hängde kvar . Men han flög ända till basen och levererade meddelandet så att trupperna räddades . 
Det var duvans förtjänst . 
Fransmännen belönade den med en tapperhetsmedalj . 
För duvor har värderingar . 
Lojalitet . Tapperhet . Integritet . 
Jag vill att ni begraver stridsyxan , i brist på bättre uttryck . 
Poängen i berättelsen är att man får ta smällar och ta på sig skulden för den stora helhetens skull . 
Ni måste vara mina Cher Ami , för jag orkar inte med fler rackarspel som det i morse . 
Ingen vill se den där Liverpool-nissen sparka in ytterdörren med sin armé av gudfruktiga vettvillingar . 
Jag förklarade för mr Dixon att jag skulle gottgöra honom om han åkte hem . 
Så nu , Eddie , måste du gottgöra mig . 
Sätt er , för fan . 
Det är som att handskas med småbarn . 
Jag har funderat igenom situationen och kommit fram till att jag har gjort mitt . 
Jack kommer att klara sig , men jag tar det som ett tecken . En uppenbarelse . Därför ska jag sälja verksamheten . 
Så enkelt är det . 
Vår överenskommelse , då ? 
Jag vill dra mig ur . Jag vill inte gå från gräsodling till massproduktion av metamfetamin . 
Jag förstår det och står fast vid det jag har sagt . Okej ? 
Inser du att du spelar mr Johnston i händerna ? 
Mr Johnston har inte en jävla susning om situationens nyanser . 
Jag tänker inte skänka bort nåt , särskilt inte till jänkaren . 
Jag tänker sälja till högstbjudande och godtar bud på 150 miljoner eller mer . Alla bud ska vara inne den här veckan . 
Jag vill att du samarbetar med Susie för att få fram den bästa dealen . 
Varför just jag ? 
Det har inte gått obemärkt förbi att ni har blivit lite av ett radarpar . 
Varför sa du inget ? 
Du har drivit verksamheten i åratal . Ska du bara låta honom sälja det ? 
Jag är bara anställd . Precis som du . 
Lägg av . Han är din pappa . Han frågade dig inte ens . 
Han frågade inte dig heller . 
Du gick bakom ryggen på mig . Två gånger . 
Vi har båda gjort en del felbedömningar , men så är det i affärer . 
Du fick som du ville till slut . 
Pappa ska sälja . Du kan dra dig ur . 
Du , då ? 
Du är för ung för att gå i pension . 
Det finns värre saker än att få sova ut och spela bingo på onsdagar . 
Ja . 
Han har bestämt sig . Det är bara att få det överstökat . 
Det är ingen hemlighet att jag vill ta över verksamheten . 
Jag är medveten om att den har stött på allvarliga störningar de senaste månaderna . 
Varor försvinner . Rutter blockeras . Smällar utdelas . 
Vi vet att du låg bakom det . Du gick över gränsen med min bror . 
Du avvisade mitt första anbud . 
Jag ville visa dig och din far att jag menade allvar . 
Jag är beredd att förhandla om ett fredligt övertagande , men du ska ha klart för dig att jag har trumf på hand . 
Ms Glass , du verkar inte känna till att en missnöjd medarbetare har försett mig med adresserna till de andra odlingarna . 
Nej , tyvärr . 
Listan mr Stevens fick var förfalskad . 
- Hallå ? 
- God dag . 
Talar jag med markisen av Beaversbrook ? 
Det är jag . 
- Baron Noughton ? 
- Hej . 
Viscount Bowling ? 
Det är jag . 
Jisses . Det här är faktiskt roligt . 
Vänta . 
Jag ringer för att diskutera er affärsrelation med mr Robert Glass . 
Ja ja . Vem talar jag med ? 
- Jag trodde att den hade kontrollerats . 
Du har blivit förd bakom ljuset , mr Johnston . 
Ja , det förvånade mig att ni två kom tillsammans . 
Varför ändrade du dig ? Det var utslagsgivande . Så jag fällde utslaget . 
Varför skulle jag vara intresserad ? 
Du har etablerade kontakter i Sydamerika . 
De skulle få en vertikalt integrerad verksamhet som har hälften av den brittiska marknaden . 
Om och när det legaliseras i Storbritannien har du en av Västeuropas mest avancerade utvecklingsanläggningar . 
Hjälpa dig ? Jag kan ordna ett möte med ryssarna , men de är jävligt råbarkade . Drar man ett skämt de inte förstår åker man ut genom fönstret . 
Frågan är om de har finanserna . 
Några hundra är en spott i havet för dem . De har Kreml i ryggen . 
Ni vet att jag menar allvar . Det har ni sett med egna ögon . 
Mina kontakter är på en annan nivå . 
Vi är beredda att ta risken . 
Och det som hände mellan oss ... 
Det bästa som nånsin har hänt mig . 
Man vet ingenting innan nån bankat skiten ur en . 
När man inser att makt är det enda som betyder nåt , öppnas världen för en . Det är bara att ta för sig . 
Din machiavelliska taktik till trots är pappa beredd att sälja verksamheten till dig , men bara om du betalar mer än alla andra . 
Förklarar det fågelns närvaro ? 
Pappa är gammaldags vad gäller affärskommunikation . 
Alla bud ska vara skriftliga och levereras med brevduvor den här veckan . 
Räcker inte ett telefonsamtal ? 
Du får fråga Bobby när du lagt det vinnande budet . 
Adjö . 
Jag älskar fågeln , förresten . Hysteriskt jävla roligt . 
Det avslutar visst våra affärer . 
- Vi har några fåglar kvar . - Vi släpper ut dem . De hittar hem själva . 
Stackars duvor . 
Lycka till . 
Lycka till . 
Det har varit känslosamt , kapten . 
Mamma , är allt bra med Geoff ? 
Han har betett sig så konstigt . 
Tja , du vet . Han har alltid tyckt om dig . Det är nog inget att bry sig om . 
Titta , där är Eddie ! 
Hej . God morgon . 
Om du letar efter din duva , så stack Freddy iväg med den förut . 
Så bra . Jag får väl gå och tygla honom , då . 
Säkert att allt är bra ? Ja , mamma . Allt är bra . 
- Vartåt gick han ? 
- Ditåt . 
Kom igen , Mitch . Ät lite . 
Då blir du stor och stark . 
Vem pratar du med ? 
Va ? Ingen alls . Pratade ? Nej , jag tror inte att ... 
Ge mig fågeln . 
Bara en duva , okej ? Bara en liten duvjävel . 
Jag vet vad du tänker säga . Du har höjdare som står i kö , men jag kan också få ihop stora summor . 
Skulder räknas inte . 
Du behöver inte raljera . Jag har sett dig under de här månaderna . Jag har sett dig hantera saker och ta in alla kriminella grejer ... 
Lyssna på mig nu . Vi ska dra oss ur . 
Inga fler spel . Inga fler skulder . Det är slut nu . 
Nu förstår jag . Du är avundsjuk . Du vill röja mig ur vägen . 
Det var du som ville röja mig ur vägen . 
Okej , det ... Jag förtjänade det där . 
- Men ... - Jag tar duvan . 
Du får inte ta Mitch . 
Du är inte ämnad för det här . 
Det är ingen av oss . 
Minns du första gången vi jagade hjort med pappa ? 
Inte direkt . 
Vi smög oss på hjorten och pappa lät mig skjuta . 
Och ta mig fan , jag prickade den . 
Han var så jävla stolt . 
Men när vi kom närmare andades den fortfarande . Det gick inte . 
Du var bara ett barn . 
Du var ännu yngre . 
Pappa gav dig kniven och du skar halsen av den utan vidare . 
Det är det jag vill ha sagt . Du kanske har rätt . 
Jag kanske inte är ämnad för det här . 
Men du ... Du är fan född för det . 
Ta hand om Mitch åt mig . 
Ursäkta att jag stör , Ers nåd , men är allt bra ? 
Du ser ut att ha det lite jobbigt . 
Inte nu , Jimmy . 
Självklart . Förlåt . 
Ta fram ett utkast till en bolagsordning . Den behöver inte vara bindande , men jag behöver riktlinjer för ett konsortium för intresserade parter . 
Vi måste nog få ihop runt 200 för att ha en chans . 
Merparten ska komma från de andra 12 lorderna . 
Om de kan gå in med tio procent var är vi på god väg . 
Sen kontaktar vi våra vänner bland resandefolket . 
De gör goda förtjänster på sin import-exportverksamhet . 
Jag har velat kapa bandet med familjen Glass ett bra tag . Jag ska ta ett kliv inåt istället för utåt . 
Det borde räcka till en plats vid bordet , men det fattas ändå en del för att nå målet . 
Om allt går bra borde ni kunna få ihop 25 , plus lånet från er mamma på tio miljoner . 
Jag fick sälja alla mina aktier och mammas Monet . 
- Tack , mamma . - Det fattas ändå 15 . 
- Okej ... - Susie Glass , då ? 
Du kan inte driva företaget utan henne . 
- Hon är inte intresserad . 
- Det har jag svårt att tro . 
Vad jag förstår har hon skött ruljangsen i flera år . 
Det är invecklat . 
Det betyder att jag måste överväga ett mindre attraktivt alternativ . 
Hej , Henry . 
- En kopp te , tack . 
- Ska bli . Du ser sliten ut . 
Du borde gå till doktorn . 
Såna här skador brukar resultera i frågor som jag inte vill besvara . 
Synd att din sponsor inte kunde hitta nån sympatisk läkare åt dig . 
Jag har i och för sig hört att dina affärer med vår amerikanska vän har nått vägs ände . 
- Varsågod . - Tack . 
Du är välunderrättad . 
Jag gav Susie de 15 miljonerna rakt av och ytterligare 15 för det där med Jack , men jag vet inte om saken är utagerad . 
Vad var det du ville ? 
Du vet vad du har gjort . Det är oförlåtligt . 
Jag vill se om det går att förändra ditt öde . 
Jaså ? 
Jag kan lösa det åt dig , men det kommer att kosta ytterligare 15 . 
Dessutom måste ett par saker fixas . 
Vad hade du tänkt dig ? 
- Hur mår han ? 
- Han sover mycket . Men han mår bättre . 
Hur mår du ? 
Jag vet inte riktigt . 
Jag fokuserar på honom . 
Ni måste stå varann nära . 
Han var tio när mamma gick bort . 
Det är ett tungt ok för unga axlar . 
Det kändes aldrig som en börda . Jag älskade att ta hand om Jack . Och jag älskar verksamheten . 
Jag vet att din pappa planerar att sälja den . Du funderar säkert på dina alternativ . 
Det enda rådet jag kan ge dig är att inte lyssna på nån , särskilt inte min son och din pappa . 
Och om du vill dra nytta av många års erfarenhet , så är det mycket mer troligt att man ångrar det man inte gjorde än det man gjorde . 
Berätta . Vad är det du tror att jag inte ska göra ? 
Jag sköter alltså grovgörat . Du tar hand om lorderna , och den där JP ... 
Sköter han distributionen ? Ja . Dina 15 gör dig till aktiv delägare . 
- Tror du att Bobby går med på 200 ? 
- Det är det jag har tänkt mig . 
När affären är i hamn är han ute ur spelet . 
Farbror Stan , då ? 
Hans redovisning har tydligen sina brister . 
Din mamma var på sjukhuset . 
Du är visst full av motsägelser . 
Kanske det . 
Är det Liverpool-hjärna uppe bland molnen ? 
Man kan hävda att han bad om det . 
Vet du vad det betyder ? 
Non sine periculo . Det är släktens motto . " Inte utan fara . " 
Det fick mig att fundera . 
Inget som är värt att ha är helt riskfritt . 
Jag insåg att släkten har sysslat med det här i flera generationer . 
Bott i en djurpark , men jagat i djungeln . 
Det är inget nytt , utan snarare upprepning . 
Har du fått ihop pengarna som krävs ? 
Vi har fått ihop en ansenlig summa , men som du vet råder hård konkurrens . 
Vi vill gärna ha fler investeringar , om du är intresserad . 
Pappa börja langa på 70-talet , för nästan ett halvt sekel sen . 
Han lyckades bygga upp ett imperium . Störst i Storbritannien . 
Men om sanningen ska fram har han tappat greppet . 
Det är som gåsen som lägger guldägg . Så länge den fortsätter värpa är allt bra . 
När jag pratat om att utöka verksamheten har han inte varit intresserad . 
Och se vad vi har åstadkommit på bara några månader . 
- Gå in med 35 , bli en jämbördig partner . 
- Vill du bli min partner ? 
Men ... vi måste prata om Henry Collins . 
Han slapp undan en gång . Det händer inte igen . 
Jag förstår . 
Men vi måste ha rimliga förväntningar , åtminstone på kort sikt . 
Du måste känna dig säker om du vill peta på den björnen . 
Oerhört . 
Charlotte . 
Låt henne flyga . 
- Redo ? 
- Kör på . 
Varsågod . 
Duktig pojke . 
Är du trött ? 
Ja , gå och mumsa lite . 
Jävlar , vilken stor siffra . 
Ja , miss Charlotte ? 
Jag har funderat en del på min barndom . 
Jag insåg att du lärde mig allt jag kan . 
Alla gånger vi campade i skogen . 
Du lärde mig att göra upp eld och rida . Hur man fångar lax . 
Det var alltid du . Eller hur ? 
Jag är bara viltvårdare . 
Är du säker på det ? 
För ibland undrar jag , och det skulle förklara en del . 
Ja , hur som helst ... 
Jag ville inte att du skulle skämmas . 
Det skulle jag aldrig göra . 
Du är den mest imponerande man jag nånsin har känt . 
Nu är fyra bud lagda . 
Alla ligger över utgångspriset . Bra gjort . 
Jag ser att ni har era namn på en av lapparna . 
Det kom som en överraskning . 
Ni ska veta att jag tänker bedöma buden baserat på deras individuella fördelar . 
- Självklart . - Perfekt . 
Men vilket bud var det som vann ? 
Det är tyvärr inte fullt så enkelt . 
Det är som ni vet hård konkurrens , och vårt bud var inte det högsta . 
Så vem vann ? 
Farbror Stan . 
Jag kände mig ganska säker på att mitt bud stod sig starkt . 
Skönt att det löste sig . 
Mr Stevens ska gå till banken och ordna så att pengarna förs över till mr Glass konto . 
Han var beredd att betala extra , så mr Glass ville undersöka budet närmare . 
Jag ser att du är misstänksam , mamma . Det är helt rätt . 
Jag hade nämligen engagerat Henry Collins , vars revisor kände till var Mr Johnston begraver sina lik . 
- Tack för att du tar dig tid . - Välkommen . 
Liken , alltså hans skatteupplägg , vidarebefordrades sedan till de relevanta myndigheterna . 
Farbror Stan greps för en rad skattebrott och fick sina tillgångar frysta . Han kunde alltså inte genomföra köpet . 
Men om han är ute ur bilden ... - Då vann väl Pete Spencer-Forbes ? 
- Det sa jag till Mercy också . 
Klibbiga Pete . 
Ditt bud kom tvåa . 
Oroa dig inte . Han vann inte . - Sa du inte precis det ? 
- Jag sa så till Mercy . 
Mina kontakter är på väg hit från Bogotá . De kommer inte att godta ett nej . 
Det är svårt att få ut pengar ur Ryssland , så det finns en liten öppning för nån som dig . 
Var finns Klibbiga Pete ? 
Mercys sydamerikanska överordnade pressade henne . 
Hon åtog sig att rensa spelplanen . 
Sen tog Henry Collins hand om henne . 
Vad skönt att nån tar hand om den stackars kvinnan . 
- Åh ... - Ursäkta . - Var det inte Henry som fixade fajten ? 
- Jo . Du jobbar väl inte med honom nu ? 
Jävla Henry Collins . 
Oroa dig inte . 
Han var desperat , så jag utnyttjade honom . 
Femton mille . Som bestämt . 
Sätt dig , Henry . 
Jag sa bara att jag tänkte sälja för att få er att vakna . 
Ni köper inte verksamheten . Ni investerar i den . 
Sen kan vi utveckla den tillsammans . 
- Du ska alltså inte gå i pension . - Va ? 
Inte en chans . 
Men jag behövde veta att ni två var beredda att sticka ut hakan . 
Delat ansvar har sina fördelar . 
Och fördelarna med kontinuitet ska man inte heller glömma bort . 
Eddie , du är soldat och aristokrat , men jag ser en man som inte låter sig definieras eller begränsas av titlar . 
Vi är alltså överens . 
235 miljoner pund . 
Nu har ni ett mål . 
Du är inte gjord för att följa order . Du ska ge dem . Du ska bygga och expandera imperier . 
Jag ser ingen kapten . Jag ser en jävla general . 
Åh , det hade du inte behövt . 
Vill du göra det ? 
Är det ett önskemål ? Nej . Du behöver inte . 
Men du kanske vill . 
Som en del av din " resa " . 
Ta det lugnt med såsen . 
Oroa dig inte . Kåken är inte så hemsk när man har vant sig . 
Man får sova ut , motionera och blir sällan störd . 
Och mr Kawasakis villkorliga frigivning drogs in , så vi kommer att äta gott i minst ett år till . 
Vad fint . 
Värre kan man ha det . 
Så talar en sann gentleman . 
