Det sägs att sorgen har fem stadier . DAG 97 
Förnekelse , ilska , förhandling , depression och slutligen , accepterande . 
Men det är nog fel att tala om stadier . Det är snarare nivåer , som i ett dataspel . 
Man kan bara gå till nivå 2 när man är färdig med nivå 1 . 
En del fastnar hela tiden på en viss nivå för att det är så svårt , som Rainbow Road i Mario Kart . 
Vilken psykopat kom på nåt sånt ? 
Allt är som det ska . 
Det är ett missförstånd . 
De är säkert vanliga , normala människor , och när de återvänder reder vi ut det här . 
" Normala människor " , va ? 
" Normala människor " , Dedo ? 
De har en hemlig bunker i trädgården . 
Och deras lilla flicka sköt dig nästan . 
Med ett armborst . 
Enligt internet finkammar de skogen efter sina nästa offer . 
Carlotta , du tror väl inte på allvar att de är kannibaler ? 
Jo . 
För tre månader sen hade jag inte trott det . 
Men då hade jag inte heller trott att min terapeut fick sin man att bära rånarluva så att hon kunde låtsas att hon hade sex med en rånare . 
Eller att min bror skulle köpa en tiger som husdjur . 
Allt det hade jag inte kunnat tro . Eller att vår dotter bara skulle försvinna . 
Och jag hade absolut inte kunnat tro att min man skulle kunna ljuga mig rätt i ansiktet i tre månader . 
Ge mig din mobil . 
Varför ? 
Vad tänker du göra ? 
Ringa polisen . De kan få ut oss härifrån . 
Ingen signal . 
Perfekt . 
Ja , det är tjocka väggar . 
Kanske även klädda med bly . 
Faktiskt rätt imponerande . 
Jackpot . 
Det är faktiskt lite romantiskt . 
Du skulle bara våga . 
De är nog preppare . 
Vad är de , sa du ? 
Preppare . Folk som tror att världen ska gå under . 
Om den bara ville komma nån gång . 
Jag jobbade med en preppare förut . 
Han var en bra jobbare . Men vi kom på att han drack sin egen urin . 
Hallå ! Släpp ut oss ! 
- Carlotta . 
- Släpp ut oss ! 
Carlotta , vi kommer på en lösning . 
Det kanske finns en annan utgång . 
Jag försöker med luckan igen . 
Hon kanske inte låste den riktigt . 
Nej . Den är ordentligt låst . 
Målet är neutraliserat . 
Presidenten informeras strax . 
Det amerikanska folket ... 
Hej . Jag visste inte vad du gillade , så jag köpte kyckling teriyaki . 
Min favoriträtt . 
Men du kunde ju vara vegetarian . Så jag köpte en vegansk macka . 
Jag är inte vegetarian . 
Okej , bra . 
Den veganska mackan såg äcklig ut . 
Okej , Chris , hör på . 
Jag har varit här nere i snart två dygn . 
De flesta som försvinner hittas inom 72 timmar . Statistiskt sett betyder det att de hittar mig här inom 36 timmar . 
Det är bara en tidsfråga . 
Det bästa för alla är att du släpper mig fri . 
Säkert . 
- Jag bara släpper ut dig , va ? 
- Jag menar allvar . 
Jag ska inte säga ett ord om dig . 
Du har varit snäll . Du köpte en smörgås åt mig . 
Jag ger dig en chans . Du ger mig en chans ? 
Okej , om du vill vara sån . 
Sundersheim är inte stort . 
Hur ofta tror du att en sexig 17-åring försvinner här ? 
- Aldrig . 
- Kallade du dig själv sexig ? 
Jag tänker sitta lugnt här och äta min smörgås , och vänta på sökpatrullen . Och då säger du ... " Snälla Wanda , tala om att jag köpte en smörgås åt dig ! " Och jag säger : " Tyvärr . 
Jag är traumatiserad och han är hemsk och borde absolut åka i fängelse . " 
Där du blir utnyttjad till höger och vänster . 
Är du klar ? 
Var ska jag gå på toan ? 
- Det är ett skämt . 
- Det här är inget hotell . 
Hur kul blir det för nån av oss ? 
Vill du verkligen bära en hink bajs uppför trappan varenda dag ? 
Chris , jag ska säga en sak . 
Du kommer aldrig undan med det här . 
Du är ingen hård brottsling . 
Polisen går från hus till hus och letar . 
De är här när som helst och hittar mig , och då åker du i fängelse ! 
Du ger mig huvudvärk . 
Sluta ! 
Låt mig gå ! 
Beklagar . 
Chris ! 
Sista chansen ! 
Jag varnar dig . Chris ! 
Chris ! 
Hur bär du dig åt , Dedo ? 
Allvarligt . 
Du tar en hemsk situation och klampar in - och lyckas göra den ännu värre . 
- Okej ... Varför följde jag efter dig ? 
Jag var ju färdig med dig . 
Det var slut . 
Jag var fri . 
Du var inte mitt ansvar . 
Men sen inser jag att du gör nåt otroligt idiotiskt igen . 
Och vad gör jag ? 
Jag följer efter dig . 
Som jag alltid gör . 
Som en idiot . 
Jag kunde ha låtit dig gå ensam , och bli skjuten av ett barn med ett armborst , och slut på historien . 
Se inte på mig som en sårad utter , som om jag ska tycka synd om dig . 
Jag tycker inte synd om dig , utan om mig ! 
Gråt inte . 
Börja inte gråta ! 
Jag gråter inte . 
- Sluta ! 
- Jag försöker . 
Jag förbjöd dig att gråta . 
Jaha , vad har de här nere ? 
Torkat kött . 
Konserverad ananas . 
Jättegott ! Konserverade bönor . 
Konserverade bönor , barbecue style . 
Jag hoppas att ni har gott om doftgranar , era psykfall ! 
Oj , toppen ! Ris ! 
Var har ni tänkt koka riset , genier ? 
Var tusan har ni tänkt koka riset ? 
Ibland roar de sig också . 
Carlotta , kanske ... Okej . 
Jaha , Dedo . 
Vad var planen ? 
Fortsätta tills pengarna är slut , och hoppas att jag inte märker nåt när de börjar utmäta våra möbler ? 
Det skulle inte gå så långt . 
Varför berättade du inte att du hade mist jobbet ? 
Vi hade hittat en lösning , vi två tillsammans , som ett lag . 
Jag kunde inte , för ... För vad ? 
Nej . 
Du hade rätt . Jag borde ha berättat . Förlåt mig . - Nej . 
Vad tänkte du säga ? - Jag tänkte inte säga nåt . 
- Jo , det tänkte du . 
Du sa " för " , och det brukar komma nåt efter . 
Carlotta , glöm det . 
För vadå , Dedo ? 
För på sistone har dina raseriutbrott blivit värre . 
Raseriutbrott ? 
Jag har inga raseriutbrott ! Jaha . 
Släpp ut oss ! Era galna jävlar ! 
Kom och ät upp oss innan vi blir skämda ! 
- Okej . - Hallå ! 
Varför gör du inget ? 
- Vad ska jag göra då ? 
- Jag vet inte ! Hitta en väg ut ! 
Kom på en plan ! 
Gör nåt istället för att bara sitta där som en idiot ! 
Det ... Oj . 
- Vad är det ? 
- Ingenting . 
Ja ? 
Den här personen tänker stanna här nere väldigt länge . 
Får hon inte ha behov ? 
Visst . Absolut . 
Var inte pryd , Dedo . 
Jag är inte pryd . Tvärtom . Jag är imponerad . 
De är verkligen väl preparerade . 
Mycket noggranna . 
Hur väl preppad måste en pervers preppare vara preppad ? 
Dedo , du är äcklig . 
Okej , bli inte arg nu . 
Jag tvättade dina kläder , som hamnade i en hög med farmors gamla kläder , och hon tog med dem till klädinsamlingen . 
Så jag gick till second hand och köpte nya kläder , men vet inte din storlek . 
Så jag kom inte till smörgåsbutiken förrän efter lunchrusningen , och då var alla goda sorter slut . 
Så jag måste köpa tonfisk ... Wanda ? 
Jag står inte ut längre ! 
Jag vägrar skita i en hink ! 
Och om jag måste äta en jävla smörgås till , kommer jag att mörda nån ! 
- Jag kan inte andas ! 
- Struntar jag i . 
Förlåt . 
Förlåt . 
Jösses . Det här är äckligt . 
Du hade nästan ihjäl mig ! 
Ja , det var tanken . 
Alltså . 
Du låste in mig här . Och du stack fingret i mitt öga , din psykopat . 
Du höll på att strypa mig ! 
Du kunde stuckit ut ögat ! 
Och jag har sagt att jag avskyr tonfisk ! 
Vad tar det åt dig ? 
Jag har varit inlåst i en gammal tants källare i två veckor ! Det är vad som tar åt mig ! 
När jag kommer ut härifrån är du rökt ! 
Du anar inte hur många poddar om sanna brott jag kommer att gå in på . 
Jag ska säga att du gjorde en massa sjuka saker med mig . 
Och alla kommer att säga : " Oj , vilken sjuk typ den där Chris är . " 
Och så ger de dig öknamnet " källarpsykopaten " . 
Och tonåringar på TikTok gör videor om dig . 
Och nån gör en film om det och nån mesig typ får spela dig . Och han säger : " Hej , jag är Chris , pervot som gillar att låsa in flickor i källaren . " 
Du är elak . 
- Är jag elak ? 
- Ja ! Du är en elak person . 
Nu minns jag . Du var elak i skolan också . 
Ursäkta ? 
Du och de andra tjejerna du hängde med . 
Ni var ett gäng med elaka tjejer . 
- Det är inte sant . 
- Jo . 
Ni höll jämt på med psykologisk krigföring på sociala medier . 
" Hur få flera gilla ? " " Vem ska jag tagga ? " 
" Hur ser jag till att alla som inte blev bjudna till partyt får veta hur häftig den är ? " Flörta med killar som visste att de inte hade en chans hos dig , tillräckligt för att de ska tro för ett ögonblick att de kanske hade en chans . För att sen relegera dem till bara vänner ! 
- Är det vad du tror om mig ? - Va ? Tror jag att du är populär och attraktiv ? Ja . 
Tror jag att det ger dig social makt ? Ja , absolut . 
Oftast är du väl inte ens medveten om vad du gör . 
Jag kan inte rå för att jag är söt och populär . Du ser ! Att du beskriver dig själv som söt och populär - är själva problemet ! - Du sa det ju själv ! 
Ja , men det är annorlunda när andra säger det ! 
Man ska inte säga så om sig själv ! 
Alltså , det kommer aldrig att hända , men anta att du sa nåt snällt om mig . 
Typ : " Chris , du är väldigt ... " 
" Du har fin frisyr . " 
Jag skulle ändå aldrig säga : " Ja , jag har fin frisyr " , för jag skulle aldrig tro på det ! 
Ska det vara nåt positivt ? 
Förlåt att jag köpte tonfiskmacka . 
Chris ? 
Du har fin frisyr . 
Händerna bakom huvudet ! Ansiktena mot väggen ! 
Jag har en AR-15 . 
En enda oförsiktig rörelse , så skjuter jag . 
- Det är ett gevär . - Ansiktena mot väggen ! 
Ja . Vi står vända mot väggen . 
Jag kommer in . Om ni inte står vända mot väggen med händerna bakom huvudet ... Händerna på huvudet . 
... ser jag det som en aggressiv handling och skjuter . 
- Uppfattat ? 
- Ja . 
Förstår ni ? - Ja , ja ! 
- Ja ! Vi förstår ! 
Herregud . 
Dedo , vad är det där ? 
Ansiktet mot väggen ! 
Vi kommer i fred . 
Vilka är ni och vad gör ni på min tomt ? 
Vi ... Vi är Carlotta och Dedo Klatt . 
Förlåt intrånget . Vi söker efter vår dotter som är försvunnen . 
Hon heter Wanda . 
Måste vi neutralisera dem , mamma ? 
Raring , nej . 
Inte än . 
Nu är de dina fångar , vännen . 
- Vill du binda dem ? - Ja . Ja ? 
Varsågod . 
Ja , utmärkt . 
Det går utmärkt . 
- Nu ! - Hallå ! 
Modigt . 
Lägg ner vapnet , annars vrider jag nacken av henne . 
Jösses , Dedo . 
Ja ! - Lägg ner vapnet ! 
- Okej . 
Gör inga plötsliga ... - Dedo ! 
- Rakt på kulorna . 
- Var det bra , mamma ? - Jättebra . Otroligt . 
Du är bäst . 
Gå upp nu . Läggdags . 
Jag tar hand om resten . 
Ge mig den . 
Älskar dig . Jättemycket . 
Älskar dig . 
Okej . Vänd er om . Händerna bakom ryggen . 
Förlåt . Det var dumt gjort . 
Det kan man verkligen säga . 
Händerna bakom ryggen . 
För hårt . 
Det skär in i huden ! Ja . Ner på knä ! 
Båda två ! 
Hör på . Jag vet inte vilka ni är . 
Men jag har aldrig sett regeringsfolk som ser ut som ni . 
Jag gissar att ni tillhör nån vänstervriden , woke , naiv gerillagrupp , visst ? Försöker skapa problem för hederliga patrioter som jag , va ? 
Förmodligen för hela KNR . 
- Vi är rökta . 
- Ursäkta . 
KNR ? 
Det nya rikets barn ! 
Som om ni inte visste det . 
Vi är bara vanliga föräldrar . 
Vår dotter försvann . 
Varför ringde ni inte polisen om ni trodde att hon var här ? 
För att polisen är totalt oduglig ? 
Där är vi i alla fall överens . 
Just det . 
Man måste slå vakt om sig . Man måste skydda sin familj . 
Nog förstår du det ? Ja . Det är sant . 
Jag litar inte heller på myndigheter . 
Därför hemundervisar jag Toni . - Gör du ? 
- Ja , hon kunde avfyra ett vapen när hon var fem . Och fånga , döda och flå en kanin när hon var sex . 
Oj , duktigt . 
Du skulle säkert göra allt som krävs för att skydda din dotter ? 
Betyder det att du släpper oss ? 
Lämna oss inte här nere ! Snälla ! 
Lossa repen åtminstone ! 
Jag har cellskräck ! 
Herregud ! 
Jag har inte cellskräck , jag bara sa det . 
Bara mord och prostitution . 
Och herr Neubert tyckte att den passade för 13-åringar . 
Vi kunde väl ha fått göra Cats ? 
Det är konstigt när man tänker på det . 
Hur gammal var du ? Tolv ? 
Perfekt ålder för att spela en hora . 
Det är det sista normala jag minns . 
Vadå ? Spela seriemördare som 16-åring ? 
Nej . 
Det var sommaren innan mina föräldrar dog . 
- Kom igen . 
- Nej . 
- Kom . Snälla , snälla . - Nej . 
Kom igen . 
- Kom igen ! 
- Okej , okej . 
Nej , " wind " . 
Ja . 
Jag har en sak åt dig . 
Herregud ! 
Det är inte sant ! 
Det fanns massor på second hand . 
Girls Team . 
Fighting Beat 2 . 
Ice Twister ? 
Mothman . 
The Mothman ! 
Jag har aldrig hört talas om dem . 
Samma här , men det kostade tre euro för allihop , så ... Alltså , jag klagar inte . 
Jag ser nu säsong två av 24 för fjärde gången , och om jag tvingas se Kim Bauer möta den där pantertanten en gång till ... 
Vad jag menar är , tack . 
Jag måste prata med dig om en sak . 
Alltså ... Jag vet att din situation är väldigt komplicerad och att de Lukas jobbar åt är superfarliga , och därför kan du inte släppa mig . 
- Wanda , jag ... 
- Nej . Lyssna på mig . 
Jag har tänkt . Om vi skulle sätta dit dem ? 
Du sa att Lukas pratade om nån " storboss " . 
Jag vet inte . Han sa " King " . Men jag vet inte om det är ett namn eller ett smeknamn . 
Okej . King . 
Alltid en början . 
Anta att det var den här King som beordrade Lukas att döda den där kvinnan . 
Frågan är : Varför han gjorde det ? 
Vad försökte han dölja ? 
- Kvinnan var journalist , va ? - Ja . Hon gjorde videor på nätet eller nåt . 
Journalist . Okej . 
Journalist . 
Om man dödar en journalist är det för att hon avslöjade nåt man vill hålla hemligt . 
Såja . 
Så om vi två kommer på vad det är , kan vi gå till polisen . Skurkarna får fängelse , jag får komma hem och du är rentvådd . 
Vi är ett team . Som Jack Bauer och Tony Almeida . 
Säkert . 
Du och jag ska avslöja den organiserade brottsligheten i stan ? 
- Ja , varför inte ? 
- Wanda . 
Jag kan inte stanna här för alltid . 
Till slut flyr jag eller smugglar ut ett meddelande . 
Eller får utbrott och slår dig i skallen med tv:n . 
Och om inte det funkar , tar jag livet av mig . 
Säg inte så . 
Jag menar det . 
Vad har jag att leva för ? 
Ice Twister ? 
Eller vi kan samarbeta och komma på en plan . Så att vi båda kommer helskinnade ur det här . 
Vad har du egentligen att förlora ? 
Jag är ledsen . 
Dedo , sluta . 
Jag är ... Jag är väldigt ledsen . 
Inte bara för det här , att få oss inlåsta i en bunker hos en beväpnad högerextremist . 
Jag är också ledsen för att jag inte berättade om uppsägningen . 
Jag ... Jag skämdes så . 
När min familj behöver mig mest , sabbar jag allting . 
- Alltid . Varje gång . 
- Dedo . Carlotta , det är sant . 
Tänk efter . 
Som när Ole föddes och läkarna sa att han var döv . Jag fick genast panik och bröt ihop , och du var den som sa : " Dedo , ryck upp dig . 
Det spelar ingen roll . Vi kommer inte att älska honom mindre för det ... " 
- Ja . 
- Och du hade förstås rätt . 
Det ändrade ingenting . 
Men i den stunden var du klippan , inte jag . 
Det var likadant när Wanda försvann . 
Sen den dagen har jag känt mig så värdelös . 
Som far är det mitt jobb att ta hand om min familj . 
Att skydda min familj . 
Och vad gjorde jag ? 
Dagen Wanda försvann , var jag berusad på en fotbollsmatch . 
Och förlåt att jag tjuvlyssnade på dig i terapin . 
Jag menade inte att göra det . Jag lovar . 
Jag hörde mitt namn och visste att jag borde stänga av , men jag kunde bara inte . 
Det var som om universum sa till mig : " Dedo , lyssna noga . 
För det här är sanningen . 
Du är en idiot och du kommer att mista allt om du inte skärper till dig . " 
Dedo , du är inte en idiot . 
Det var fel av mig att säga så . 
Men du hade rätt . 
Jag är en idiot . Jag har alltid varit en idiot . 
Det var så jag drog mig fram i livet . 
Det var så jag kom genom skolan . 
Det var så jag fick dig . 
Dedo , den älskvärda idioten . 
Ingen har höga förväntningar på en idiot . 
Om man gör bort sig blir ingen förvånad . 
Man får sämre betyg och sämre lön än andra ? Det är ju sån Dedo är . 
Dedo , du tror väl inte på det där ? 
Vet du inte vad ... du betyder för mig ? 
Carlotta , varje dag är jag rädd att du ska säga : 
" Dedo , allt det här var ett misstag . Jag vill skiljas . " 
Men det händer inte , av nån anledning . 
Kanske är det för att vi fick barn så tidigt , så du kanske känner att du är fast med mig . 
Jag vet inte . 
Jag älskar dig så , Carlotta . 
Att gifta mig med dig var det bästa som nånsin hänt mig . 
Och när jag ser dig le mot mig på morgonen vill jag ropa av glädje . 
Och jag frågar mig varje morgon : 
" Dedo , hur tusan gick du i land med det här ? " 
Jag förstår det inte . 
Jag förstår inte varför nån som du står ut med en sån som jag . 
Jag förstår det inte . 
- Jag ville bara ... - Nej . 
- Var tyst . - Okej . 
Dedo , dra ner blixtlåset på mina byxor . 
- Okej . Det är en knapp också . 
Okej . 
- Känner du den ? 
- Ja . - Kan du ... 
- Ja . 
- Det går . 
- Bra . 
- Kom hit nu . - Ja . 
Okej . - Lägre ner . - Bra . 
Lite till . 
- Lite till . 
- Såja ! Åh . Herregud . 
- Okej . 
Vänta . Vänta lite . 
- Nej . Lite längre ner . - Okej . 
- Åh , jösses . - Åh , jösses . 
Åh , jösses . 
DAG 68 ... visst ser hon hemsk ut ? 
Det är nog ! Jag går hem . 
Det är nog ! 
Jag är ingen ... Sluta filma mig ! 
- Dra åt skogen , allihop ! - Herregud . 
Ledsen , Wanda . 
Jag borde inte ha visat dig videon . 
Nej , det var bra att du visade mig den . 
Jag ... Jag känner mig så skyldig . 
Blunda ett tag . 
Varför ? 
Bara blunda . 
Okej , men gör inget knäppt . 
Jag känner mig rätt skör just nu . 
Okej . 
Nu kan du titta . 
Vad är det där ? 
Jag visste att videon skulle göra dig ledsen , så jag tänkte muntra upp dig och köpa all din favoritmat . 
Nattvickning ! 
Först av allt en ananas . 
För på din allra första utlandssemester lät din pappa dig smutta på hans piña colada . 
- Och du sa att det var ... 
- Det godaste jag nånsin smakat . 
Nachos . 
Sweet chili , för du älskar hur kryddstoftet fastnar på fingrarna . 
Och oliver för du tvingade dig själv att tycka om dem , så folk skulle tycka att du var sofistikerad . 
Och sist men inte minst ... Strängost . 
Jo , och för gamla tiders skull ... Bara lugn . Det är inte tonfisk . 
Kom du ihåg allt det där ? 
Det var nog det snällaste nån har gjort för mig . 
När jag fyllde år senast fick jag en kokbok för en varmluftsfritös av min dåvarande pojkvän . 
Jag har aldrig ägt en varmluftsfritös . 
Alltså , jag menar inte att du är min pojk ... Vänta , jag har en sak till . 
- Ja ? 
- Ja . 
Jag kan inte . 
Förlåt . 
- Jag menade inte att ... 
- Det är inte så att jag inte vill . 
Det är snarare tvärtom . 
Jag menar , hallå ? 
Du är den snyggaste tjej som nånsin har pratat med mig . 
Fast det är inte det . 
Du är rolig och smart och så totalt oberörd av hela världen . 
Och jag har aldrig mött nån som är så tuff och modig som du . 
Men jag vill inte vara en läskig kille ... Och ja , jag vet att jag håller dig inlåst i min källare , - vilket är superläskigt ... 
Slappna av . Det är okej . 
Nog för att jag har tänkt på det . 
Jag är ju kille och hetero . 
Det är bara ... Vänta , titta . Jag googlade . 
" När maktbalansen är ojämn kan det vara svårt att avgöra om medgivandet är frivilligt , och genuint medgivande kan även vara omöjligt . " 
Just det . Och därför går jag min väg nu och önskar dig en trevlig kväll . 
Hej då . 
Jag har diskuterat saken med min dotter . 
Vi är båda mycket upprörda över ert olaga intrång . 
Och tyvärr är min bunker inte helt laglig , så om ni anmäler det här hamnar jag i en stor knipa . 
Vi ska inte säga nåt . Jag svär . 
Vänd er om . 
- Du behöver inte . - Vänd er om . 
Jag älskar dig . 
Och jag dig . 
Faktum är att jag förstår . 
Som en mor . 
Om Toni försvann skulle jag söka ända ner i helvetet efter henne . 
Och efter att ha gjort en snabbkoll på nätet är det tydligt att ni två inte är hemliga agenter för djupa staten . 
- Just det . Ja . - Ja . 
Dedo , du bör ompröva din närvaro på sociala medier . 
Du lägger ut många memes . 
Många . 
Och de är inte bra . 
Jag ska ta det under övervägande . 
Hoppas att ni finner henne . 
Jag vet inte vad jag skulle göra om jag miste Toni . 
Bara så att allt är klart : Är vi fria att gå ? 
- Ja . 
- Okej , då går vi . 
Jag lämnar den här . 
Jo , vi drack lite av din vodka . 
Och jag åt upp en burk lasagne . 
Jag vill gärna ersätta den . Dedo . 
Om du ger mig dina bankuppgifter - kan jag över ... - Mm . 
Tack så mycket för din förståelse . 
Oss mödrar emellan uppskattar jag det verkligen . 
En sak till . 
Det är ett litet hål i ditt staket . 
- Jag kan ... 
- Dedo . 
Det är inte sant . 
Vem är du ? 
Tack för titten , morfar . 
Wanda . 
Farmor gav mig just det här . 
INSATSGRUPP WANDA KLATT En polis var här och frågade om min skåpbil . 
En insatsgrupp bara för mig ? 
Coolt . 
Vadå ? 
Det här kanske är nåt bra . 
Om de vet om din skåpbil , kanske de vet om Lenka och Lukas också ? 
De letar inte efter Lukas , utan efter mig ! 
Lugna ner dig . 
Det ordnar sig . Vi löser det här . 
Tillsammans . 
Vi måste sluta . 
Sluta att spionera och göra intrång och ljuga för polisen . 
Men jag menar inte att vi ska ge upp . 
Vi fortsätter leta . Men inte så här . 
Vi måste vara rädda om det vi ännu har . 
Ta hand om oss själva och Ole . 
Annars finns inget kvar för Wanda att komma hem till . 
DAG 97 Presidenten informeras strax . 
Det amerikanska folket ... Ojsan . 
Farmor ? Det är Chris . 
Är allt bra ? 
Plötsligt slocknade lyset . 
Oroa dig inte , jag kommer hem nu . 
Nej , det behövs inte . 
Jag har ringt Lukas . 
- Lukas ? - Okej , jag ska ta en titt . 
Var är säkringsskåpet ? 
I farfars gamla hobbyrum . 
Är det nån där ? 
Hallå ? 
Är det nån där ? 
Chris ? 
Wanda . 
- Vi måste härifrån . 
Är det nån där ? 
- Kom nu ! 
- Vänta . 
Vad gör du ? 
Wanda , kom nu ! 
