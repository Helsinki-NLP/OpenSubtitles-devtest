Denna serie är ett fiktivt verk . Den är inspirerad av historiska händelser , men platser , personer , organisationer och händelser i detta drama är fiktiva . Tidigare i Uncle Samsik 
Angående herr Choo ... 
Beordrade du hans mord ? 
Du låter fantasin flöda igen . 
Varför visa honom Innovationspartiet ? 
Han var besatt av nationalförsamlingen ... 
Förbered eldgivning ! 
... så jag trodde att en nominering skulle tysta honom . 
För att hedra min far måste vi skingra oss omedelbart . 
Det ska inte utövas nåt mer våld . 
Ser du ? Inget hände . 
Det vet vi inte än . 
- Var är Cha Taemin ? 
Jag hittade Sineuialliansens uppförandekod , signerad av Kang Seongmin , men Pak Jiwook brände den . 
Signerad av Kang Seongmin ? 
Men han brände den ? 
Jag erkänner att jag var med i Sineuialliansen . Jag formulerade deras uppförandekod . 
Svär du på att du inte dödade min son ? 
Yoon Palbong och jag dödade An Minchul i Cha Taemins ställe eftersom han förrådde Kang Seongmin . 
Ge mig en chans . 
En sista chans . 
Jag övervakar dig . 
Kang Seongmin vill få igenom lagen om lokalt självstyre . 
Det är din chans att etablera din närvaro . 
Ska jag gå emot honom ? 
Vi vill få igenom lagförslaget så att han kan avancera i Liberala partiet . 
Lagförslaget är ogiltigt ! 
Jag har inget mer att lära dig . 
Genom att motsätta mig framstår jag som en kämpe för demokratin . 
Det är nåt skumt med Samsik . 
Han har umgåtts med Kim San , Choo Intaes svärson . 
Vem är Kim San ? 
- Du ska få ett större scoop . 
- Ett scoop ? 
En bild värd förstasidan på bråk i Nationalförsamlingen . 
Bra jobbat . 
Jag gör det . 
Militären kan försöka ge förste infanterichefen makten . 
Första infanterichefen ? 
General Choi Hanrim . Militären litar på honom och han står nära USA:s befälhavare . 
Du är väl bekant med general Choi ? 
General Choi passar perfekt som vår affärspartner . 
Du bör ansluta dig till oss . 
Jag planerar en statskupp . 
Vi behöver logistikkommandots hjälp för att flytta trupper och utrustning snabbt och diskret . 
Vi börjar förbereda när datumet är satt . 
Jag tog in general Choi . 
Och jag valde dig . 
Välj mig , så följer familjen Albright med . 
Du verkar ha turen på din sida . 
Vi ska stjäla hans perfekta plan . 
Vad är din plan ? 
Jag tar Pak Jiwook med Han Soo som lockbete . 
Och sen ? 
Sen tar jag Choi Hanrim med Pak Jiwook . 
Jag ska stoppa hans dröm om en statskupp . 
Jang Doosik blir befälhavare för kapitalförsvarsenheten och Jeong Hanmin vice befälhavare . 
Då hamnar Choi Hanrim i Jang Doosiks och Jeong Hanmins våld . 
Från och med idag är du Kim Kwangmin , Sanaekoncernens vd . 
Vi bad om att få betalt i mjöl för exporten av råmaterial i enlighet med givarlandets begäran . Och vi vill få mjölet till den officiella växelkursen . 
" Då får ni mer än fem gånger så mycket betalt . " 
- De bygger en bro åt dig . - Vi bygger en bro . 
Jag föreslår att de får mjölet till den officiella växelkursen . 
Då får Sanaekoncernen betalat enligt den officiella växelkursen ? 
Vi har aldrig setts , okej ? 
Vad var det i den där lådan ? 
Kang Jinseong ? 
- Kang Seongmin . 
Sineuialliansens stadgar . 
Pak Jiwook måste ha gömt dem . 
- Varför skulle han göra det ? 
- Pak Jiwook måste planera ... - Ja ? ... att hugga Kang Seongmin i ryggen . 
Pak Jiwook ... 
Uncle Samsik 
Uncle Samsik 
Tvivel 
- Han är här . - Han är här . 
Erkänner du anklagelserna ? Kommentera . 
En kommentar , herrn ? 
Åklagarna har bevis på att du tog emot mutor . 
- Ur vägen . - Sluta . 
Vem har tutat i er det ? 
Avgå , Pak Jiwook ! 
Lugna ner er , allihop . 
Liberalernas ledamot Pak Jiwook anklagas för mutbrott 
Okej . 
Han är på Nationalförsamlingen . 
Okej . Jag tar en påtår . 
Kaffet är extra gott i dag . 
Har du lagt till nåt speciellt ? 
Kärlek och omtanke , såklart . 
Det är därför det smakar så gott i dag . 
Nationalförsamlingen 
Gjorde du Sanaekoncernen en tjänst gällande deras exportintäkter ? 
Nej . 
Varför den officiella växelkursen ? 
Det var kommitténs kollektiva beslut . 
Du visste att de skulle få mer än fem gånger marknadsvärdet , va ? 
Alla i kommittén var överens om det . Skyll inte på mig ! 
Vad är det med er ? 
10 mars 1960 Seoul , Sydkorea Hotell Banya 
Vart är Korea på väg ? Av journalist Choo Yeojin 
Val påverkade av regeringsmanipulation , mutor ... 
Varje tecken på korrupt demokrati uppenbaras framför våra ögon . 
Med maskopi , konspiration och skenhelighet verkar valet bli än mer förvirrat . 
Vi får se om detta politiska kaos blir Koreas växtvärk eller dödsdom . 
Prova den . 
Vad är det ? 
En kostym till dig . 
Vad tycker du ? 
Du ser bra ut . 
Svär eden . 
Jag ser dåligt . 
" Under dagens utfrågning ... " 
" Under dagens utfrågning ... " " ... som hålls av Nationalförsamlingen i mutfallet ... " 
" ... som hålls av Nationalförsamlingen ... " 
Från och med i dag är du Kim Kwangmin , Sanaekoncernens vd . 
- Välkommen . 
- Här borta . 
Hej . Jag är Kim Kwangmin , vd för Sanaekoncernen . 
Han ser för ung ut . 
Han är äldre än han ser ut . 
- Berätta vad du behöver . 
- Ja . 
Vi bad om att få betalt i mjöl för exporten av råmaterial i enlighet med givarlandets begäran . Och vi vill få mjölet till den officiella växelkursen . 
- Du kan hjälpa oss . 
- Va ? 
När vi får betalt i mjöl ... 
Det betyder att ni får mer än fem gånger så mycket betalt . 
Du har rätt . De ger dig 20 % av vinsten och en bro i din valkrets . Vad säger du ? - En bro ? 
- Ja . 
- Kan han göra det ? 
- Givetvis . 
Jag gör allt du ber om . 
Jag gör mitt bästa . 
Lägg det diskret i bakluckan . 
Ja , herrn . 
Hej då ! 
Vilka är ni ? 
Varför står ni i vägen ? 
Vi är från åklagarmyndigheten . 
Åklagarmyndigheten ? 
Och ni har fräckheten att stå i vägen för en ledamot ? 
Ta honom . 
- Håll fast honom . - Släpp ! 
Släpp , sa jag ! 
Bad ledamot Pak dig om valfinansieringen först ? 
Ja , han behövde pengar . 
Sa han det själv ? 
Ja . 
Så du erkänner anklagelserna ? 
Vad betyder det ? 
Mutade du honom ? 
Ja . 
Tala klarspråk . 
Jag mutade honom . 
Pak Jiwook går inte fri . 
Vittnena vittnade mot honom . 
Är Sanaes vd Kim Kwangmin ett vittne ? 
Känner du honom ? 
Han är Kim Sans vän . 
Här kommer han . 
Demokraterna för ekonomin ! - Choo Intae ! - Choo Intae ! - Choo Intae ! 
- Demokraterna vinner ! 
Var han vittnet ? 
Han är inte Kim Kwangmin . 
Vittnena blev förväxlade . 
- Leverera det här . 
- Va ? - Förväxlade vittnen ? - Ja . 
Gå och berätta för dem . 
Det är till dig . 
Säger du att vi förväxlade vittnena ? 
Va ? Ett falskt vittnesmål ? 
Var är vittnet nu ? 
- Vittnet . - Ja ? 
Är du medlem i Dongdaemunligan ? 
Ja . 
- Gav du falskt vittnesmål ? 
- Ja . 
Så du vill ändra ditt vittnesmål ? 
Ja . 
Men du försåg ledamot Pak med politiska medel ? 
Ja , det stämmer . 
Det var min chefs order . 
Känner ni till Yoon Palbong ? 
Han sköts till döds av Sineuialliansen . 
Så du gav de politiska medlen till ledamot Pak på Yoon Palbongs order ? 
Ja , precis . 
Vad var anledningen ? 
Ingen aning . Jag följde bara order . 
Sluta med det där . 
Så du följde hans order ? 
Det är mitt jobb att följa order . 
En fråga till . 
Träffade du ledamot Pak genom Daemyeon Byggs vd Yoo Yeonchul ? 
Vem är det ? 
- Din jävel ! - Herrn . 
- Vem är du ? 
- Sa du jävel ? 
- Vem fick dig att göra detta ? - Säg det igen ! Han saknar hyfs . 
Yoon Palbong beordrade mig att vinna över ledamot Pak . 
Mutan kom från honom . 
Varför gjorde Yoon Palbong det ? 
- Hur ska jag veta ? - Varför inte ? 
Jag vet inte . Jag ... 
Jag menar ... Jag följde bara min chefs order . 
Nånting stämmer inte . 
Vad menar du ? 
Jag presenterade Yoon Palbong för min far . 
Det är ett nöje . 
Jag heter Yoon Palbong . 
Kände du Yoon Palbong ? 
Jag kommer strax . 
Vart ska du ? 
Kan jag hjälpa dig ? 
Vilken organisation tillhör du ? 
Vad är kopplingen mellan Jiwook och Kwangmin ? 
Kände du Yoon Palbong från Dongdaemunligan ? 
Ja . 
Kim Kwangmin presenterade honom för Innovationspartiet och kontaktade mig med flit . Sen sköts Yoon Palbong tillsammans med min far . 
Har det inget med min far att göra ? 
När träffade du Kim Kwangmin ? I går . 
Vi borde inte prata här . 
Vi pratar nån annanstans . 
Jag vet inte var jag ska börja , men Pak Jiwook satte dit flera oskyldiga medborgare under japanskt styre . 
Herr Choo var en av dem . 
Om han har satt dit andra , är det väl rätt att sätta dit honom ? 
Jag menade inte så . 
Varför gick han med i Innovationspartiet ? 
Han ville väl bli ledamot . 
Vem övertalade honom ? 
Det kan jag tyvärr inte berätta . 
Så du vet . 
Nån försöker döda Pak Jiwook och Yoon Palbong . 
Det är allt jag vet och allt jag kan dela med dig . 
Kan jag tro dig ? 
Ja . 
Våga inte bråka med min far . 
- Släpp . Kang Seongmin . 
- Lugna dig , herrn ! 
Släpp . 
Vi måste prata . 
- Journalisterna hör dig . 
- Det struntar jag i . - Kang Seongmin . 
- Övertygade Yoon Palbong dig ? 
Va ? 
Jag undrar vems order han lydde . 
Misstänker du mig ? 
Utfrågningen kommer nog att klargöra allt . 
Du , Kang Seongmin . Du kan inte göra så här . 
Du borde inte ha gjort så här . Vad har jag gjort ? 
Sineuialliansens uppförandekod . 
Du hade bränt den . Men du ljög . 
Du borde ha förvarat den på ett säkert ställe , inte åkt runt med den i bakluckan . 
Här , herrn . 
Hej . 
Kan du få det gjort i dag ? 
Jag måste se det innan jag svarar . 
Det måste ske inom en dag . 
Om du lyckas dubblar vi summan . 
Då ska jag göra mitt bästa . 
Den här vägen . 
- Varsågod . 
- Okej . 
Sineuialliansens uppförandekod " Sineuialliansen ... " 
Vad är det här ? 
Bry dig inte om vad som står . 
Hur fort kan du göra en kopia ? 
Tja ... 
Räcker det om jag är klar vid midnatt ? 
Tar det så lång tid ? 
Du behöver bara skriva några bokstäver . 
Det är inte ... så enkelt . 
Håll det hemligt . Om du är klar inom tre timmar betalar vi mer . 
- Mer ? 
- Ja . 
Det här också ? 
Okej . 
Vem ? 
Choo Yeojin ? 
Träffade du henne igen ? 
Drog du in herr Choo ? 
Jag är upptagen . Låt mig ... 
Varför sa du inget ? 
Lägg inte på nu . 
Du borde inte träffa henne igen . 
Hon kom hit . Hon varnade ... Hon varnade mig för att bråka med hennes far . 
Okej , jag tar hand om det . 
Hur då ? 
Jag kommer över . 
- Är det kampanjschemat ? 
Det är många som vill höra ditt tal . 
Bra jobbat . 
Kan du skilja dem åt ? 
- Inte alls . 
- Vilken är originalet ? 
Kan du inte knacka eller nåt ? 
Vad gör du ? 
Jag försöker ruinera Kang Seongmin . 
Vilket är originalet ? 
Det här ? Det vänstra ? 
Vilket är originalet ? 
Det till vänster . 
Då är det denna . 
Snygg kostym . 
Kan vi prata lite ? 
Ny kostym ? 
Var är Kwangmin nu ? 
Han är i Nationalförsamlingen . 
Presenterade han Yoon Palbong för Yeojin med flit ? 
Vad gäller det ? 
Svara mig . 
Ja . 
Vd Kim är här . 
Var fick du kostymen ? 
Byt inte ämne . 
Nån har bra smak . 
Använde du Kwangmin också ? 
Varför gjorde du så mot herr Choo ? 
Bara få general Choi att lämna militären . 
Du bryr dig om Choo Yeojin . 
Det är inte poängen . 
Vem köpte kostymen ? 
Svara nu . 
Var det Rachael ? 
Blåsfisken ? 
Vill du inte svara ? 
Vill hon att du deltar i statskuppen ? 
Vill du delta ? 
Nej . 
Jag tänker sätta dit Choo Intae tillsammans med Choi Hanrim för spionage under Arbetarpartiets 29:e direktiv . 
Varför sa du inget ? 
Det dök nyss upp . 
På Kang Seongmins order ? Ja . 
Du bryr dig om honom . 
Sanaekoncernen fick betalt i mjöl för deras exportintäkter . Du gjorde orättvisa vinster genom den officiella växelkursen . 
Jag blev förvånad över betalningen . 
Bad inte du ledamot Pak om en tjänst ? 
En logistikofficer nämnde hans namn . 
En logistikofficer ? 
Vem ? 
Kapten Kim Inho från kapitalförsvaret . 
Varför träffade du logistikofficerarna ? 
Jag gör affärer med armén . 
Vad sa kapten Kim ? 
Att Yoon Palbong bett om en tjänst . 
Vad för tjänst ? 
Att presenteras för högt uppsatta militärer och politiker . 
Vilka politiker syftar du på ? 
Nämn bara namnet Pak Jiwook vid förhöret . 
Jag lovar att du inte råkar illa ut . 
För ett hederligt liv behövde du släppa din girighet . Men du ville ha både lutfabriken och Cheongwooförbundet . 
Man får bara tillfredsställa några begär . 
Ingen får alla . 
Det är givet . Så vad ska vi göra ? 
Du borde öka dina begär . 
Har du inga ambitioner ? 
Han nämnde ledamot Pak . 
Vilket skitsnack ! 
Vem är du ? 
Samsik ligger bakom det här , va ? 
Din jävel . 
Jag blir ditsatt ! 
Det är en lögn ! 
- Släpp ! 
- Det här blir rörigt . 
Vilken huvudvärk . 
Vem är Kim Inho ? 
Kära nån . 
Ursäkta mig . 
Du utreds av CIC , eller hur ? 
- Ja , herrn . - På vilka grunder ? 
I relation till Arbetarpartiets 29:e direktiv . 
Utveckla vad det är . 
Det hänvisar till Nordkoreas spionage för att vinna över vår militärpersonal . 
Varför var en medlem i Dongdaemunligan inblandad i spionaget ? 
Yoon Palbong lydde visst under Nordkorea . 
Yoon Palbong ? 
Han som sköts av Sineuialliansen ? 
Ja , herrn . 
Jag hörde att han fick order på kortvågsradio och levererade en taltabell för att dechiffrera dem . 
Till vem ? 
Kapten Pak Wonil från kapitalförsvarsenheten . 
Det är gåvor , herrn . 
Gåvor ? 
Jag beställde dessa åt dig från en affärsman som importerade varor till logistikkommandot . 
Jag har redan mutat kapitalförsvaret . Hong Youngki har planterat bevis med Arbetarpartiets 29:e direktiv . 
Du ville väl ha en bok ? 
Ja , ordnar du det ? 
Den kan skickas från Japan . 
Tack . 
Gillar du Choo Intae ? 
Du , det går att vinna . 
Hur då ? 
Den avlidne Choo Intae . 
Ska vi använda en död person ? 
Vi använder honom eftersom han är död . 
Samexistensens stig 
Vad står på ? 
Min far är deras mål . 
Var Samsik inblandad i mordet på Choo Intae ? 
Nej . 
Det var en olycka . 
Menar du att Choo Intaes död var en olycka ? 
Pak Jiwook var ditt lockbete . 
Du visste allt , va ? 
Ska du döda general Choi med hjälp av Pak Jiwook ? 
Ja . 
Allt föll på plats . 
Varför gömde du general Choi ? 
För att utnyttja honom bakom ryggen på Samsik ? 
Du planerade det med Jeong Hanmin och ordnade ett gömställe åt general Choi . 
Hej . 
Välkommen . 
Hur gick det ? 
Jag har en plats åt general Choi . 
Tack , Hanmin . 
Jag visar dig en annan utgång . 
Jag möter dig där . 
Lystring ! 
President Rhee kommer att vara i sitt fritidshus på valdagen . 
Stället vaktas av runt 20 personer . Den 122:a bataljonen är stationerad i närheten och består av 500 soldater . 
Den 15 mars , dagen för presidentvalet , är vår bästa chans . 
Var redo att offra era liv för ert land ! 
En dödspatrull på 30 man från armén , tusen från logistikkommandot , femhundra från 55:e Howitzerregementet , och 1 000 från 31:a divisionen kontrollerar Jinhaes semesterhus . Kapitalförsvaret och 3:e marinkårsregementet blockerar vägarna till huvudstaden . 
Vi tar radiostationer , Bank of Korea och tågstationer i storstäderna och utfärdar order om undantagstillstånd . 
Kapitalförsvarskommandot 
Vi hittade den i din vas . 
Förklara . 
03 attack , 04 påbörjas , 05 hemligt möte 
Okej . 
Min Soochul har gripits . 
Vi borde återgå till våra baser . 
Vi borde nog det . 
Herrn . 
Vi borde skynda oss till baserna . 
Du kan inte åka tillbaka . 
Va ? 
Du kommer att gripas så fort du kommer dit . 
Jag eskorterar dig till en säker plats . 
Följ med mig . 
Vi är nästan framme . 
Kim San . Vad gör du här ? 
Jag eskorterar dig härifrån . 
Följ mig . 
Herrn . 
Var är general Choi ? 
Gick inte han ut tidigare ? 
Hur gick det ? 
Vi missade general Choi . 
Vad pratar du om ? 
Han var vårt mål ! 
Hur kan du dricka nu ? 
Jag njuter inte av det . 
Letar dina män efter Choi Hanrim ? 
Jag undrar hur han fick reda på vår plan . 
Nån kanske har gömt honom . 
Vet du vem som ligger bakom ? 
Varför gömde du general Choi ? 
Var du verkligen inte med på statskuppen ? 
Vi vet inte var general Choi är än . 
Vi säger till så fort vi vet . 
Får du tag på Kim San ? 
Nej , det får jag inte . 
Märkte du inget misstänkt ? 
Skulle jag ha märkt nåt misstänkt ? 
- Varför gör ni så ? 
- För bort dem ! 
- Vänta ! 
- Släpp mig ! 
Vad pågår här ? 
För bort henne . 
Ni har ingen rätt att storma ett partikontor ! 
Vad gör ni ? 
För att dechiffrera nordkoreanska sändningar använde de Choo Intaes böcker , inklusive Fredlig återförening och Samexistensens stig . 
Under Arbetarpartiets 29:e direktiv , försökte spionen Choo Intae vinna över flera högt uppsatta politiker och militärer . 
Han verkar också ha etablerat Innovationspartiet för att utföra uppdraget . 
Du gör mig galen . 
Har du kollat upp Yeojin ? 
Jag vet inget . 
Lägg av , okej ? 
Hon kan väl släppas ? 
Jag vet inte , sa jag . 
Vad är det med dig ? 
Tack , herrn . 
Choo Intae visar sig vara nordkoreansk spion 
Hur länge måste jag vara här ? 
Tills presidentvalet är över . 
Det dröjer inte länge . 
Vad händer där ute ? 
Vi undersöker det . 
Planerade ni att gömma mig här i förväg ? 
Ja , herrn . 
Varför då ? 
Choi Minkyu ville bli av med dig och använda dig i valet . 
Jag fick information från inrikesministeriet . 
Choi Minkyu ? 
Du har rätt . Det är effektivt . 
Den allmänna opinionen har vänt . 
Utländsk media förväntar sig ett jämnt val . 
Vi kan vända på situationen . 
Jag har en idé . 
Låt mig komma över . 
Nej , jag kommer över . 
Det visade sig vara effektivt . 
Klyftan mellan de två partierna minskade snabbt . 
I hur många regioner leder Demokraterna ? 
Det finns 20 regioner där de leder stort . 
Klyftan är för stor . 
Vi kan inte vinna här med legitima åtgärder . 
Föreslår du att vi ingriper på nåt sätt ? 
Vi måste stjäla valurnorna . 
Herrn , det är ... 
Det går bra om vi vinner . 
Om vi vinner får vårt agerande nu inga konsekvenser . 
Hur ska vi stjäla alla valurnor ? 
Samsik sköter det . 
Det är hans specialitet . 
Jag behöver tänka lite . 
Det hinner vi inte . Valet är nära . 
Ring honom nu . 
Ska jag ringa ? 
Sineuialliansens uppförandekod Kang Seongmin 
Det här är min signatur . 
Du har räddat mig igen . 
Jag har haft svårt att sova på grund av det här . 
Du kan sova gott nu . 
Tror du att jag kan bli premiärminister ? 
Självklart . 
Du är nästan där , herrn . 
Choi Minkyu har ännu ett orimligt krav . 
Vadå ? 
Men det är inte rätt . 
Berätta för mig . 
Vi ligger långt efter i vissa regioner . 
Säg inte att du vill ha valurnorna ... 
För riskabelt ? 
Jag menar ... Jag har stulit allt möjligt , men aldrig valurnor . 
Okej . 
Glöm att jag nämnde det . 
Situationen kommer väl inte att vända ? 
Det blir ett jämnt val , men vi leder i stora områden . 
Ser ni ? Vi leder stort i alla områden där Kim San kampanjade . 
Du blir säkert nominerad . 
Jag vill bara ha nationell rekonstruktion . 
Kom igen . 
Bekymra dig inte för det . 
- Ursäkta mig . - Okej . 
Vad gör du här ? 
Saken är den ... De har gripit Yeojin . 
Va ? 
De kanske inte släpper henne . 
Kan du hjälpa till ? 
Vad tittar du på ? 
Du borde ha sagt att du var här . 
Det gjorde jag . Vad tittar du på , sa jag . 
Det är inget . 
Låt mig se . 
Kang Seongmin bad mig ... 
" Valdistrikt där demokraterna leder " ... stjäla valurnorna . 
Är han galen ? 
Choi Minkyu fick honom att göra det . 
Försvarar du honom ? 
Vad pratar du om ? 
- Nu är du löjlig . 
- Tänker du stjäla dem ? 
Nej , jag ska få honom att glömma det . 
Lura inte dig själv . 
Vissa saker kan jag inte förklara . 
Jag har inga såna . 
- Är du säker ? 
- Ja . 
Gav Rachael dig nåt annat än kostymen ? 
Vad ska det betyda ? 
Hon erbjöd nog en position efter statskuppen . 
Jobbar du på reformen åt mig ? 
Vad gör du här så här sent ? 
Polisen har gripit Yeojin . 
Kan du få ut henne ? 
Då blir det komplicerat . 
Så du vill inte . 
Det sa jag inte . 
Bryr du dig så mycket om henne ? 
Ja . 
Hon kommer att stå i vägen för oss . 
Okej då . Strunta i det . 
Jag kan göra det . 
Men det blir bara jobbigt . 
Ska du stjäla valurnorna ? 
Jag ska få ut henne . 
Är du nöjd nu ? 
Menar du att du slöt ett avtal med Samsik på grund av Choo Yeojin ? 
