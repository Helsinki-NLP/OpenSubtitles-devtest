Hörru , grabben ! 
- Får han låna skrivbordet ? 
- Javisst . Slå dig ner . 
Vet du hur illa det här är ? 
Jag har en viss aning . 
Jag kan fixa undan kroppen , om du vill ha hjälp med det . 
- Han , då ? 
- Herr Tvångssyndrom som räknar pengar . 
- Vi kan ta hand om honom också . 
- Vi kan inte döda honom . 
- Har du nåt bättre förslag ? 
Fyra miljoner prick ! 
Knäpptyst . 
Jag fattar . 
Han får skylla sig själv . 
Kom hit ! 
Jethro ! 
Stanna , för fan ! 
Hej , Geoff . 
- Vad är det vi jagar ? 
- En blå träningsoverall . 
Freddy , kör norra vägen . 
Jag går österut . 
- Vet du vart du ska ? - Jadå . 
Ingen mottagning ! 
Stanna , Jethro ! 
Hämta andan , grabben . 
- Det räcker . 
- Jag ska inte säga nåt . 
Jag såg inget . Okej ? 
- Gör mig inte illa . - Det ska vi inte . 
- Vi löser det här . 
- Va ? Ni dödade ju Tommy ! 
Jag lovar . Vi ska inte göra dig illa . 
Okej . Nu avslutar vi det här . 
Lägg ner vapnet . 
Inga vittnen . 
Vad fan är det med dig ? Ge hit den där . 
Släpp mobilen . 
Släpp mobilen , Jethro . 
Freddy , nej ... 
Mobilen är rökt . Bra där . Nu kan du berätta vem han skulle kontakta . 
Låt dem komma . 
Låt de jävlarna komma . 
Kom nu . 
Vad fan betyder det här ? 
Vi lider alla med dig , Johnny . 
Vi vet varför du är här . 
Du har övergett dig själv i den fysiska känslans vildmarker . 
Det handlar inte om bilen eller klockan på din handled . 
Det handlar inte om de fem grammen koks eller vad han nu tar på fredagskvällar . 
Du vet att den marken är ofruktbar . 
Därför är du här . Därför är vi alla här . 
Vi kan erbjuda dig ... kärlek och broderskap . Världen där ute kan inte erbjuda dig nåt förutom en kista full av ihåliga ben . 
Så slut ögonen och öppna ditt hjärta för Gud . 
Okej , då tar vi en stund för att reflektera . 
Maxie . Ta över . 
Ursäkta , John , men vi får inte tag i Tommy . 
- Han svarar inte i telefon . - Och ? 
Han skulle hämta pengarna . Nu är han borta . Han hittar väl på nåt bus . 
Jag brukar inte oroa mig , men jag fick ett sms från Jethro . 
Vad stod det ? 
Det var tvetydigt . 
Vad menar du ? Otydligt . Öppet för tolkning . 
Jag vet vad tvetydigt betyder , Errol . Vad skrev han ? 
Okej . Vi måste förvara honom nånstans tills det här är utrett . 
- Hur stor är din frys ? 
- Inte stor nog . 
- Går det att låsa arbetsrummet ? - Ja . 
Stäng fönsterluckorna , lås dörrarna . Ingen går in . 
- Hur många finns i huset ? 
- Mamma och 20 anställda . 
Ge personalen ledigt resten av dagen . Sen avvaktar du . 
Tjugo anställda , ledigt . Uppfattat . 
- Edward , ha koll på honom . - Ja . Överlåt det åt mig . 
Kom , då . 
Du . Bilen . Nu . 
Okej , sätt dig . 
Prata bara med personalen , ingen annan . Det är lugnt . Lugna puckar . 
Det är bara mycket att smälta . 
Det känns som om allt är i 3D . 
Allt är i 3D . 
- Ja , men det känns annorlunda på nåt sätt . 
- Det är annorlunda . För du har mördat nån . 
Ska jag bara stå här och titta på honom ? 
Får jag göra mitt jobb ? Gå på toa ? 
Jag vill att du aktiverar skallen , Jimmy . 
Vad i helvete ? 
Jag vet inte om det går . Jag behöver tydliga instruktioner . 
Det går bra . Det är bara några timmar . 
Låt honom inte använda telefonen . 
Han är vår fånge och i knipa . 
- Låt honom inte snacka sig ur det . 
- Okej , chefen . 
Inga problem . 
Röker du gräs ? 
Hur så ? Har du nåt ? 
Vi måste lösa det här utan att fler blir dödade . 
Det sista nån av oss vill ha är fler lik . 
Det är rörigt . Och dåligt för affärerna . 
Men du måste förstå vad vi har att göra med . 
Tommy Dixon var ganska långt ner i näringskedjan . Men hans bror , Gospel ... Han är lite mer att bita i . 
Och en jävla blådåre . 
Han är farlig . Och han känner mäktiga personer . Vilka då ? 
Jesus . Och hans farsa . De har gjort honom till en av de största kokainlangarna i nordväst . 
Jesus och hans farsa ... Tuff kombo . 
Förliten eder icke på furstar , icke på en människoson . Han kan icke hjälpa . 
Hans ande måste sin väg . Han återvänder till den jord varav han är kommen . Då varda hans anslag om intet ! 
" Jag är vägen , sanningen och livet . Ingen kommer till Fadern utom genom mig ! " 
Vedergällningen manifesterad . 
Du behöver inte vara med . Låt oss proffs sköta det . 
- God morgon . - Bonjour . 
- Felix , är allt bra ? 
- Utmärkt , tack . 
Jag skulle precis kliva upp , faktiskt . 
Jag har ett jobb åt dig . 
Har du tid idag ? 
Idag ? 
Jag ska kolla min kalender . 
Du har tur . - Men nån måste köra . 
Jag måste ... Dra igenom listan igen . 
Kalk . 
Fluorvätesyra . 
- Vad är det ? - Bensåg . 
- Såg ... - Sticksåg . Stickande såg . 
- Plastpåsar . - Påsar . 
- Och skyddsdräkter . - Va ? Skydds ... 
Då kör vi . 
Och vi behöver kaf ... fe . 
Kaffe . 
Hur började du med det här ? 
Jag var med i kyrkokören . 
Jag gillar musik och siffror . 
Det är det musik är , siffror som rör sig i samklang . 
De erbjöd mig jobbet . Att sköta räkenskaperna . 
Jag visste inte att de var en gangsterfamilj . 
Tommy Dixon framstod inte som särskilt religiös . 
Där tar du fel . 
Den här Jesusförgreningen är dödligare än senapsgas . 
Bröderna är helt från vettet . 
Det enda de gillar mer än kärlek är att mörda . 
Tommy förtjänade det . 
Skönt att han är död . 
Jag ska inte säga nåt . Jag svär vid Jesus . 
Den andra Jesus . Den snälla . 
Jag kanske tror dig , men det är fler som ska övertygas . 
- De kommer att döda mig . 
- Inte nödvändigtvis . 
Upp och hoppa , Felix . 
Felix . Buongiorno . Du ser ut att vara i form . 
Blanket , kan du öppna bakluckan och ta fram mattan ? 
Det fixar jag . 
Det är kallt . 
Då så . Är läget under kontroll ? 
I nuläget . Mamman sover där uppe . Personalen har fått ledigt . 
Okej . Ett lik och ett vittne , va ? 
Inga konstigheter . Är vittnet säkrat ? 
Då börjar vi med liket . 
Vad fan väntar ni på ? 
Om ni ska med får ni klä av er . 
Okej . Ett kadaver med en svår huvudskada . 
- Är det där vapnet som användes ? 
Är det en Gainsborough ? 
Fantastiskt . 
Vi får putsa den sen . 
Det får bli ett kapa och gräva-jobb . 
Vi delar kroppen i fyra delar , letar reda på en fridfull , avskild plats , begraver den djupt , strör över kalk , packar gropen med jord och dekorerar med gödsel . 
- Jag har en fråga . 
- Varsågod . Varför måste den delas ? 
Då kan man gräva ett mindre hål . 
Och när de inre organen exponeras , påskyndar man förmultningen . 
Maskarna älskar det . 
I mitt yrke måste man tänka holistiskt . 
Keith , tvätta bort blodet från väggarna . 
Blanket , lägg vapnet i bilens bagageutrymme . Ställ bilen på baksidan , så att den är utom synhåll . 
Jag styckar kroppen där ute . 
Utför du operationen ? 
Ja . Jag erbjuder full service , inklusive undanröjandet av vittnen . 
- Fler frågor ? 
Då kan vi hälsa på värden . 
Eddie , det här är Felix . 
Han har gott om erfarenhet av såna här situationer . 
- Han erbjuder sin expertis . 
- Hej . Hej . Tack för att du kom så snabbt . 
Ja , tiden är ju av vikt . 
Jag uppskattar din expertkunskap , men vi måste prata om Jethro . 
Är Jethro vittnet ? 
Vi kan utnyttja honom för att skapa en alternativ historia för Gospel . 
Jag kan antyda att nåt var på tok mellan Tommy och Jethro . De tjafsade medan han räknade pengarna . 
Vi filmar uppträdandet med Tommys mobil . Sen lägger vi kroppen i bilens baklucka . 
Då tror Gospel att Jethro dödade Tommy och tog pengarna . 
Ursäkta , men var är Jethro när allt det utspelar sig ? 
På ett fraktfartyg till Australien . Med två mille i fickan . 
Det vore enklare att skicka honom till Lappland . 
Han kan chilla med tomten , gömma sig bland nissarna och bygga leksaker . 
Det är en bra kille som råkat i trubbel . 
Han behöver bara få andra alternativ . 
Vad tycker du , Felix ? 
Ni borde hugga huvudet av honom . 
- Toppen . - Jag vet vad din pappa skulle göra . 
Han skulle också hugga huvudet av honom . 
Lyckligtvis sitter han inne , så vi slipper . 
Utmärkt . Då var det klargjort . Håll kvar Jethro , så pratar jag med Gospel . 
Städa huset , men gör dig inte av med kroppen . 
- Ursäktar du oss lite ? 
- Visst . 
- Vi går och pratar . - Gärna det . 
Du verkar ha glömt varför vi är här . 
Jag försöker hjälpa dig att lösa problemet . 
Om du inte vill ha min hjälp ber jag Felix packa ihop . 
Nej . Jag ber om ursäkt . 
Jag vill inte verka otacksam . Jag behöver bara lite tid för att se om jag kan lösa det här . 
Mord är dåligt för affärerna , sa du . 
Tjugofyra timmar . Sen måste vi städa . 
Bra . 
Jag vill inte göra det . 
Jag ville inte förut heller . 
Jag tänker fan i mig inte dansa . 
Du gjorde nåt väldigt dumt , Freddy . 
Du dödade nån . Det kan inte göras ogjort , men om du gör exakt som jag säger finns det en liten chans att du kommer undan med det . 
Du ska dansa . 
Okej , då . 
Mr J. 
Använder ni Waterman Serenity-bläcket ? Blått , inte svart ? 
Det stämmer . 
Se till att använda läskpapper . 
Jag vill lägga till ett namn på gästlistan . 
Skicka en inbjudan till hertigen av Halstead . Se om han nappar . 
Så där . 
Jag är en sprätt som tabbade mig Lian , lian , lej 
- Bäst hittills . 
- Ja , men ändå dåligt . 
- Nämen , älskling ... 
- Hej , mamma . - Vi ska bara göra en grej . Behöver du nåt ? 
- Det här levererades precis med bud . - Okej . 
- En inbjudan från mr Johnston . 
Johnston med ett " T " ? 
Ja . Känner du honom ? 
Inte formellt sett . 
Vad synd att det inte var du som fick inbjudan , då . 
Vill era vänner ha te ? Ja ? Personalen är som bortblåst . 
Te vore gott . 
Jag kan ta hand om det . 
Tack , Geoff . 
Det är nog på tiden att jag träffar Stanley Johnston . 
Jag trodde att vi var klara med honom . 
Lapsang souchong . 
En kaka ? Tack , Geoffrey . Vad snällt . 
Frederick , varför är du klädd som en höna ? 
Ja , precis . 
Alltså , hönan är lite av en ... Grejen med hönan är ... Vad skulle du säga , Eddie ? 
- Välgörenhet . - Just det . Välgörenhet . 
För vadå ? 
En organisation som uppmärksammar de hemska förhållandena för burhöns . 
Exakt . Vad altruistiskt av dig . 
Jag visste inte att du brydde dig om djurens väl och ve . 
Man gör det man kan , för hönsens skull . 
Jag är lite förvirrad , ms Glass , men vad exakt är det du jobbar med ? 
Min man sa nåt om antikviteter , men nu verkar du så engagerad i djurens välbefinnande . 
Vilket är det ? Antikviteter eller höns ? 
Jag har inget intresse för bristerna inom kommersiell hönshållning . 
Hans nåd har välsignats med ett mer medkännande hjärta . 
Jag har hjälpt honom med affärerna och ville stötta honom . 
Skål för det . 
Nu har han ringt tre jävla gånger . 
- Tror du att han vill prata med mig ? 
- Det får man nog anta , ja . 
Om det här ska funka måste du bete dig som om allt är bra . 
Okej , jag vill inte vara taskig , men grejen är att du måste svara . 
- Hallå . Freddys mobil . - Är Freddy där ? Jag vill tala med honom . 
Tyvärr inte . Ska jag hälsa honom nåt ? 
Jag heter John Dixon . 
Vem pratar jag med ? 
- Edward , hans bror . 
- Okej . Ett sånt sammanträffande . Det gäller nämligen min bror , Tommy Dixon . 
- Har du hört talas om honom ? 
- Ja , han var faktiskt här i morse . 
Just det . Det är bra att veta . 
Han har inte kommit hem , så jag undrar var han är . 
Han åkte härifrån runt kl. 11.00 . 
- Och du var där ? 
- Ja . 
Då är du den sista som har sett honom . 
Det var tråkigt att höra , mr Dixon . 
Kan vi hjälpa till på nåt sätt ? 
Kan jag titta förbi imorgon vid tolvtiden ? Då kan vi prata igenom allt . 
- Javisst . Om det är till hjälp . - Det är det . 
Då så . Ta hand om dig till dess . 
Errol , det luktar trubbel . 
Imorgon klockan tolv ? Bravo . 
Freddy , varför kommer det två bilar ? 
- De tog med hela gänget . 
- Ingen lätt packning här . 
Låt er inte skrämmas av mina killar . 
Det är bra killar . Gudfruktiga . 
God dag , mr Dixon . 
Är det din kåk ? Ja . 
Väldigt ... Versace . 
Imponerande . 
Driftkostnaden måste vara chockerande . 
Vad är det för nåt ? 
- Du känner visst min bror , Freddy . 
- Ja , vi känner varann . 
Du borde göra bot . För Jesus älskar dig . 
Vi känner varann väl . Så bra . 
Mr Lawrence . 
Varsågoda . Ta med hela kören . 
Vad tråkigt att höra att din bror är försvunnen . 
Som jag sa i telefon : När Freddy var klar igår morse , åkte de . Vi har inte hört nåt mer . 
Löstes affären till Tommys belåtenhet ? 
Dra åt helvete ! 
Ja . Freddy gav Tommy pengarna . Tommy väntade medan hjälpredan ... 
Jethro , va ? 
- Ja . - Ja . Jethro kontrollräknade pengarna och sen gav de sig av . 
Problemet är att ingen av dem har hörts av sen de åkte härifrån . 
Sen fick vi ett kryptiskt sms från Jethro . 
Errol , visa dem meddelandet . 
" Tackla Tommy Woo Woo . " 
Är det nåt religiöst ? Det tror jag knappast . 
Nej . Kan han ha haft mobilen i fickan ? 
Kanske det . Men jag tror att han ville ha nåt sagt . 
Frågan är ... vad . 
- Eddie , har du nån aning ? 
- Nej , tyvärr . 
Men det var en sak ... 
Det är nog inget , men det inträffade en mindre dispyt . 
Vad menar du ? 
- Det är när två ... 
- Jag vet vad det betyder . 
Medan Jethro räknade pengarna blev din bror frustrerad . Det blev en ordväxling . 
- Låter det likt dem ? 
- Jag har aldrig hört dem vara osams . 
Vad var de oense om ? 
Tommy blev frustrerad över att det tog sån tid . Jethro ville inte ha nåt tjat . 
Tommy är inte den mest tålmodiga . 
Det kanske inte var mer än så . Det kanske inte var nåt . Precis . Jag hopps att Tommy bara har avvikit från vägen . 
Det vore inte första gången . 
Det finns inget Gud älskar mer än en syndare som återvänder till fållan . 
På tal om det , är det nån här som behöver göra bot ? 
Är det nåt du vill berätta , Frederick ? 
Ja . Jag har en bekännelse . 
Jag har tagit ett liv . 
Vem har du dödat ? 
Förlåt , Eddie . 
Jag bar ansvaret för Montys död . 
- Katten Monty ? - Ja . Nån sa att man kan lära en katt simma genom att kasta den i en sjö . Så jag kastade i honom . Han åkte i plurret och sjönk . 
Jag letade efter honom i två veckor . Förlåt . Det var 25 år sen . 
Jag trodde att det var en trygg zon . 
Nåt mer ? 
Ja , jag pullade den där hushållerskan som du gillade ... Freddy . 
Vad fan gör han ? 
Tack för att ni tog er tid . Ursäkta att jag störde . 
Ingen fara . 
Hoppas att du hittar honom . 
Tack . Men jag tror inte det längre . 
När jag stod där borta fick jag en överväldigande känsla av att min brors själ har lämnat hans kropp . 
Jisses . 
Det är storartat på sitt sätt ... För att visa respekt vill jag hålla en tyst minut . 
Går det bra ? 
Ja . Absolut . 
- Ska du ... - Edward , kan du ... 
Vill du ... 
Vi borde nog ... 
Oj , vilket hårt grepp . 
Hell dig , Maria . Amen . 
Okej , nu drar vi ! 
Köpte han det ? Det känns så . Det är nog för tidigt att avgöra . 
Ja . 
Om han gjorde det , om vi tar oss igenom det här , ska jag gottgöra dig . Jag pratar inte om pengar . - Då är jag skyldig dig mitt liv . 
- Ja , det är du . 
Lägenhet 12 , sjätte våningen . Passet ligger i strumplådan . Tredje lådan , bakom kallingarna . 
Och du delar inte lägenhet med nån ? 
Jag bor ensam . 
Okej . Jag fixar det . 
Vilken hektisk dag . Så mycket folk . 
- Väntar vi fler ? 
- Nej . Det var nog allihop . 
Jag vet att det är svårt att ha folk springande här , men det är inte för alltid . 
Vad skrattar du åt ? 
Din pappa sa nåt liknande . 
- Tack , Lawrence . 
- Ers nåd . 
Men det fanns inget han kunde göra åt det . 
Du visste . - Ja . - Du har vetat hela tiden . 
Varför sa du inget ? 
För att du måste fatta ett eget beslut . 
Din pappa såg inga fel med det . 
Pengarna gagnade oss alla . Men det förgiftade honom . Det förgiftade hans själ . - Jag vill inte se det hända dig . 
- Det ska jag inte tillåta . 
Men nu måste jag hantera en sak . - Freddy ? - Ja . Freddy . 
Men när det är gjort ska verksamheten bort från godset . 
Okej , men ... lova att vara försiktig . 
Om man lämnar en glipa i luckan smyger sig naturen in . 
De blir väl förvirrade . Det är som permasommar här nere . 
Det kommer allt möjligt . Snokar , hermeliner ... 
En gång flög en rödhake in . 
Jag fångade den som en baseboll . 
Vet du att om man lägger pekfingret på rödhakens huvud och juckar som mellan två tuttar och får till rytmen helt rätt , så ger fågeln sig till en . 
Benen särade , vingarna åt sidan . 
Det är jag . - Hej . - Säg att det inte är där han sa . 
Han säger att det han letar efter inte är där det skulle vara . 
Det trodde jag . 
- Han säger att det är där . 
- Va ? - Kollade han strumplådan ? 
- I lådan . - Jimmy . - I lådan . Ge honom telefonen . 
Jag har strikta instruktioner om att inte ge honom nån telefon . 
För då kan han ringa nån . Och han är ju vår fånge . 
Fråga igen var passhelvetet är . 
- Det ska ligga i strumplådan . Vänta . - Fan . - Det ligger under keyboarden . - Va ? Spelar du keyboard ? - Han spelar keyboard ! - Jimmy ... - Jag är rätt bra . 
- Jag har också spelat . - Jimmy . - Kolla vid keyboarden . 
- Under den . 
- I ett skåp . - I ett skåp . 
- Jag vet inte vilket , men det är litet . - Okej . 
Fan också . 
God kväll . 
Tack . 
Ser man på . Klädd som en krigare . 
Fixade du passet ? 
Gick det bra ? 
Du ser sliten ut . 
Vad gör vi här ? 
Vi undrar varför farbror Stan erbjuder mer än godset är värt . 
Varför säger du " vi " ? 
Det är nog inte huset han vill ha , utan vår verksamhet . 
- Har han en egen ? - Meth . Har tjänat miljarder på det . 
Och vad är du ? 
En knarklangare med hjärta ? 
Vi gillar pengar lika mycket som alla andra . Men hans grejer har ett våldsamt pris . 
Vi håller oss till vår relativt fridfulla marknad . 
Släpper vi in honom , blir det blodbad . 
Där är ni ju . 
Mr Johnston är mån om att få ert sällskap . 
Varsågoda . 
Hans nåd , hertigen av Halstead , i sällskap med sin vän , ms Susie Glass . - Välkommen . - Ursäkta dröjsmålet . 
Jag sprang på en vän . Angenämt . 
Tillåt mig att presentera prinsessan Rosanne . 
- Hej , Rosie . 
- Eddie . 
Rosie , Eddie , Ers nåd , Ers Höghet ... 
Vi tillbringade somrarna på Halstead förr . 
Det var länge sen . 
Det borde jag ha anat . Världen är liten . 
Prinsessan Rosanne är ättling till kung Leopold III . - Hon är elva i den belgiska tronföljden . 
- Tolva , trodde jag . 
- Vem har vi förlorat ? 
- Pappa föll av hästen . Beklaga inte . 
Du gillade honom inte . 
Han hade sina förtjänster . Den främsta är du . 
- Vad tråkigt med din pappa . 
- Verkligen . 
- Kände ni hertigen ? 
- Susie arbetade med honom i åratal . 
- Inom vilket fält ? - Jag är antikhandlare . 
Ett sånt sammanträffande . 
Då kanske ni kan reda ut en sak åt oss . 
Jag passar på att prata med prinsessan medan ni polerar antikviteter . 
God kväll . 
Din bror kan inte vara glad över att bli förbigången . 
Det har varit en utmaning . 
Har svaret varit koks och partajande ? 
Mycket av det förstnämnda , mindre av det andra . Ursäkta . Det här är mrs Jones . 
Det här är Susan Glass . 
Så trevligt . 
Mrs Jones ger mig råd om förvärv . 
Hur känner du mr Johnston ? 
Han är väldigt underhållande och generös . 
Jag har nyligen köpt en speciell klocka . 
Mrs Jones har bett mig göra en kopia . Nu undrar jag om ni kan se skillnaden . 
Jag noterade att det är en Patek Philippe 1518 . 
Så observant av er , ms Glass . Det är inte bara det . 
Det är klockan Winston Churchill bar när han accepterade Tysklands kapitulation 1945 . 
- Vet du vad han jobbar med ? 
- Vad det än är så gör han det bra . 
Han skickar jämt privatplan , presenter och yachter ... 
Jag förstår . 
Vad säger du , Susie ? Hur mycket är den värd ? 
En Patek Philippe från den tiden brukar gå för 2,5-3,5 miljoner , men med tanke på historien , att den var med när fredsavtalet undertecknades , skulle jag säga mellan nio och tio miljoner . 
Tio poäng . 
Just därför insisterade jag på en kopia . 
- Och vad får han av dig ? 
- Han får umgås med en prinsessa . 
Du har säkert märkt att han samlar på aristokrater . 
Ms Glass , kan ni berätta om klockan är äkta eller falsk ? 
Om du vill vara så snäll . 
Den är äkta . 
Förargar det dig att han bär den ? 
Det gick fort . Hur kan du veta ? 
En kopia skulle kännas varm . 
Äkta kristall är svalt tack vare lägre konduktivitet . 
Eller så chansade jag bara . 
Jag köper inte kopior . I min värld behöver jag inte det . 
Ens rykte kan lösa alla säkerhetsproblem . 
Om jag lämnar klockan på bardisken vet jag att den ligger kvar när jag kommer tillbaka . 
Det ger oss tid att röka en cigarr . 
Ska vi gå ? 
Hoppas att du vet vad du ger dig in i . 
Han är en riktig gentleman . 
Vet du vad du ger dig in på ? 
Så pinsamt . 
Jag läcker visst . 
Ska vi snygga till dig ? 
Ja . 
- Så där . - Tack . 
Ska vi sätta igång , ms Glass ? 
Låt oss inte låtsas att vi är som de . 
De lever i en djurpark , medan vi lever i djungeln . 
Berätta då varför du sniffar runt i min del av skogen . 
Din pappa har gjort ett enastående jobb med att göra verksamheten lönsam . 
Och du har varit duktig på att undvika konflikter och konkurrens . 
Men den formeln håller inte längre . 
Varför inte ? 
Om det ändå vore som förr . 
Du behöver en partner . 
Är du ett jävla orakel , eller ? 
Vad tror du att du vet som jag inte vet ? 
Du har helt rätt . 
Jag ser framtiden . 
Och om du vill att saker ska förbli som de är , så måste nåt förändras . 
Tja , tack för visat intresse . Jag ska fundera på saken . 
Ring inte mig . Jag ringer dig . På vägen ut ... - Glöm inte gåvan . - Gåvan ? 
Klockan . Den är till dig . 
Klockor får man när man går i pension . 
Din tajming är fel . 
Fan . Försiktigt . 
Stå still . 
Kapten . 
Hej , Susan . Är allt som det ska ? 
Vi täpper till ett hål . 
Klart . 
- Vad har du gjort med honom ? 
- Tja , det ser ut som en skottskada . 
- Vad har du gjort med honom ? 
- Dumma pojke . 
Det hände nog inte här . 
- Jag vet inte om jag vill veta . 
- Det vill du nog inte . 
Edward , ring mig . 
Jag hittade passet , men priset var lite högre än förväntat . 
Välkommen till djungeln . 
Måste jag ringa Felix ? 
Redan gjort . 
Vad betyder det ? 
Han är på plats med strikta instruktioner . 
Ska vi sätta igång ? 
Tack , Felix . 
Det här är planen . 
Lyssna noga . 
När Gospel ringer döingen ... 
- Döingen ? - Ja . Döingen . Det här är din värld , inte min . 
- Det var självförsvar . 
- Ta det lugnt . 
När Gospel kommer och letar hittar han kroppen . 
Varför det ? 
Vi lämnar den där . Som om Jethro dödade honom när han letade efter sitt pass . 
Gospel kommer att förstå allt när han hittar Tommy och hagelgeväret i bakluckan på bilen vid båtkajen . 
Så ironiskt . Du skulle rädda en mans liv och dödade en annan . 
Ironin går inte obemärkt förbi . Ser jag ut att behöva läxas upp ? 
Det är ingen uppläxning , utan en observation . 
Ska vi dra ? Tänker du hjälpa en gammal soldat ? Eller bara stå där och hytta med fingret ? 
Det går bra . 
Sätt dig , så tar jag av dig skorna . 
Här . Ta ett järn . 
- Klarar du dig ? 
- Ja , med det här . 
Är du kvar ? 
Inbilla dig inget . 
Jag ligger inte med personalen . 
Natti natti , mördaren . 
Vem ska nu ta av mig skorna ? 
Vänta här . 
Sändaren i hans Merca gav ifrån sig ett livstecken . 
Vi hittade den parkerad vid lotsbåtskajen vid Themsen . 
Det här är en kista , inte en bil . 
Den här låg i hans ficka . Bevisföremål A. 
På den finns videon med din brors ursäkt . 
Så det verkar som om ni hade rätt . 
Där har vi den . Det var inget helhjärtat uppträdande , va ? 
... kuk-kuk där ... Säg inte det . 
Det krävdes faktiskt en del ansträngning . 
Jag är en sprätt som ... Jethro visade sig vara en riktig vessla . 
Hur då ? 
Han mördade två män och försvann med pengarna ! 
- Har ni hittat honom ? 
- Det kommer vi att göra . Var så säker . 
Det är bara en sak som bekymrar mig . 
Vapnet min bror sköts med låg i bilens baklucka intill liket . 
Skjutvapen eller kniv ? 
Det är ett finare engelsktillverkat jaktgevär . 
Det är tydligen värt över 200 000 pund . 
Hur fick Jethro tag i det ? 
Det finns en enkel förklaring . Geväret är mitt . Eller vårt , åtminstone . Det var pappas . 
Jag märkte att det var borta när ni hade åkt . 
Vapenskåpet står ofta olåst , slarvigt nog , och ingen hade koll på Jethro . 
Jag tänkte väl att det var ert . Det är inte direkt förstavalet för en langare från Liverpools bakgator . 
Det här är dess naturliga miljö . Det var därför jag tog med det . 
Jag ville återföra handen till handsken , så att säga . 
Men på vägen hit utvecklades en utomvärldslig kontakt mellan mig och den där yttersta domens doning . 
Det kanske är mycket begärt , men kan jag få behålla geväret ett tag ? 
- Det kan bli knepigt rent juridiskt . 
- Då kan vi råka i klistret . 
- Men ... - Eller så behåller du det . 
Så vänligt . 
Var så säkra : Domen kommer att uppenbara sig . 
Och då återlämnas geväret . 
- Vi får nog tacka Jesus för det där . - Amen . 
Kan vi återgå till det lugna livet nu ? 
När du pratar om det lugna livet ... Undrade du aldrig var pengarna kom ifrån ? 
Vet inte . Slaveri ? 
Jag måste visa dig nåt . 
Jävlar i min lilla låda . 
Välkommen till djungeln . 
Den där båten tar dig till ett fraktfartyg mot Australien . 
Det är som ett tåg som stannar överallt , så det tar tid , men det är säkrast så . 
Vad var det du försökte skriva i meddelandet till Gospel ? 
" De dödade Tommy , SOS . " 
- Hur blev det " woo woo " ? 
- Prediktiv text , antar jag . 
Det är svårt att skriva när man jagas genom skogen av arga hundar . 
Lycka till . Tack . 
- Honom ser vi inte igen . 
- Du har säkert rätt . 
Du , jag uppskattar hjälpen , men den ursprungliga överenskommelsen gjordes mellan våra fäder . 
Det är dags att jag träffar honom . 
Det kan ordnas . Bra . 
Är det nåt jag kan ta med ? 
- Han älskar att grilla . 
- I fängelset ? 
Det är en öppen anstalt . 
Och han har vissa privilegier . 
Det är en fantastisk filé . 
Underbar marmorering . 
Och vilka vackra ryggbiffar . 
Verkligen . Det var vänligt , Ers nåd . 
Georgie , öppnar du taket ? 
Du måste ha bra kontakter . 
Pappa hade parkboskap på ägorna . 
De är kommersiellt ohållbara , men de håller vandrare borta . 
Stora horn . Taskig attityd . 
Jag gillade din pappa . Det var en bra man . 
Du kan gå , George . 
- Jag är tillbaka till solnedgången , då . 
- När är jag nånsin sen ? - Va ? Du är jämt sen , för fan ! - Stick iväg med dig . 
Jag sparar en köttbit till dig . 
Vet ni varför det heter " sirloin " ? 
På 1600-talet hade kung James , en avlägsen släkting till dig , en bjudning med över 100 rätter . 
I slutet av den andra dagen serverades han en bit kött som var så jävla mört och smakrikt att han dubbade den till riddare . 
" Res dig , sir Loin . " 
Begreppet fastnade . 
Och resten är historia . 
Fan , ursäkta . Sätt dig , för guds skull . 
Sätt fötterna under bordet . Värm knäna . 
Tack . 
Inget slår en grillning mitt i vintern . 
Jag måste erkänna att det här inte var vad jag väntade mig . 
Det här är inget . 
Vi har en golfbana med nio hål , en nordisk bastu och en damm vi kan bada i . Gör underverk för cirkulationen . 
- Men är inte knivarna ett problem ? 
Fängelsedirektören är en beundrare av mr Kawasakis prisade hantverk , som vi strax ska få avnjuta . 
Var det nåt du ville fråga mig ? 
Går det bra ? 
- Inför honom ? - Ja . Du kan prata öppet . Mr Kawasaki är pålitlig . 
Om det inte gäller att betala skatt . 
Eller hur , kocken ? 
Ärligt talat är det oklart om det gagnar mig att ha verksamheten på min mark . 
Jag skulle vilja öppna för nya förhandlingar . 
Vänta lite nu . Ursäkta mig ? Går vi inte händelserna i förväg nu ? 
Det skulle vara en förutsättningslös träff . 
Lite spott på fingrarna innan du matar bävern . Vi skulle inte omförhandla nåt . 
Din pappa verkar vilja höra vad jag har att säga . 
Vad har du tänkt dig ? 
Jag vill att ni försvinner före årsskiftet . 
I gengäld garanterar jag att ni tjänar mycket mer pengar . 
Mr Kawasaki , lägg biffen på grillen . 
Och häll upp lite japansk whisky åt oss . 
Vi ska visst ha ett riktigt möte . 
Du borde ha tagit upp det med mig först . 
- Du klampade över gränsen . - Du hade vägrat . Klart som fan . 
Du är en soldat ur adeln , inte en knarklangare från södra London . 
Vänta . Det var jag som sa det . Du behöver mig för att sluta döda folk . 
Vi gillar inte att döda folk . Vem fan gör det ? 
Det var din kokainsniffande bror som satte oss i klistret . 
När man väl börjar döda , måste man slutföra det . 
Jethro , då ? 
Han får gå , va ? 
Han är ju redan borta . 
Det är kallt ute . 
Kom in hit . 
- Ja , gärna . Tack . - Ja . 
Värm dig med en kopp te . 
