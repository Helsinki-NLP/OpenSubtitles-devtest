Kära vänner , det är här vi äntligen anländer till vår stora vandrings hjärta och själ . 
Det här är Market Street ! 
Men mycket har förändrats sedan jag ägde ett hus i korsningen av Fourth . Men en sak är sig lik : Unga Ava säljer brownies så mäktiga att kung George skulle försöka beskatta dem , utan laga kraft . 
Så ge er ut , goda medborgare , och spendera era pengar ! 
Som alltid är du dagens höjdpunkt , Benji . Åh , efterrätt ! Kan jag få en blondie ? 
Tryffelbrownien är min favorit . 
Känner jag igen dig från någonstans ? 
Kanske från frimurarlogen ? 
Nej , jag menar allvar . 
Har du varit i Kansas City ? 
Jag tror inte det . 
Är det ett av koloniernas nya distrikt ? 
Unga fröken , vet du vad mer som hände här på Market Street ? 
Jag gjorde mitt berömda experiment med elektricitet . 
- Titta vad jag hittade , morfar ! - Jag får se . 
Oj , den är fin . 
Avundsjuk ? Nej . 
Skojar du ? Jason får lov att ha vänner . Jag vill inte kolla Waynes bakgrund . Jag ber bara om en tjänst . Jag förstår det , men ... 
Vänta . Visst var det rummet tomt ? Har du anställt någon ? Nej . 
- God morgon . - God morgon . 
Rosa till Batista . - Och lila till Adebayo . 
- Kemi går bra . - Ursäkta , vem är du ? 
Helen , er nya kriminaltekniker . 
- Jag har inte begärt mer personal . 
- Inspektör Braun har skickat mig . - Har han placerat dig här ? 
- Jag trodde att han hade sagt det . 
Överraskning ! Jag älskar överrask - ningar - särskilt de med gåvor . 
Varsågoda , öppna dem . 
Jag börjar . Se där . 
Åh , presenter ! 
- Åh , är det ... 
- Ett krämägg från Cadbury . 
De är så goda . 
Jag fattade inte riktigt , men Cadbury är aldrig fel . 
- De är jättegoda . 
Tack så mycket . - Trevligt att träffas , Helen . 
- Jag måste ringa inspektören . 
- Ni glömde den här ! 
- Jag ser fram emot att jobba här . - Okej . 
Om du inte stannar för att köpa kaffe , måste du ta med kaffe . 
- Det var inte jag som var sen . 
- Du ville att vi skulle köra ihop . 
Ja , för Braun kommer att hålla koll på oss . 
Jaha , är du min barnvakt nu , eller ? 
Nej . Jag är din partner . Om du inte beter dig som ett barn . 
Okej , partner . 
Jag har tänkt mycket på Maritz bilbomb . 
- Snälla , låt bli . 
Maritz kommer ut och sedan smäller det . 
Undrar du inte ? Jo , men jag tänker på Nikki . Braun var tydlig . Fallet tillhör mordroteln . 
Försvåra inte för henne med den nya chefen . Var professionell , släpp det . 
- Ska jag vara professionell ? - Ja . 
Professionell som i att sjunga om en förlovning inför hela kontoret ? 
- Jag sjöng häcken av mig . 
- Det är inte poängen . 
Jag stämde av med HR . Det var ett vackert ögonblick . 
Ja , ett vackert , oprofessionellt ögonblick . 
Om du säger det så . 
Hej , Kemi . 
Skönt att du ringde , för Mike skulle precis sjunga för mig . Ska du också fria till honom ? Vad trevligt . 
Ser du ? 
Oprofessionellt . 
Erkänn bara ! 
Är ni i närheten ? 
Vi har en märklig situation här . 
- " Benjamin Franklin " saknas ? 
- Jag kan inte ljuga . Vår nations grundare och landsman har försvunnit . 
Vi jobbar som historiska vandringsguider . 
Jag heter Alexander Hamilton . 
Vissa av oss är strikta med att inte gå ur sin roll . 
Det menar ni inte . 
Franklin försvann under en rundtur i dag , men var alltid ett proffs . Mer inne i sin roll än George . 
Han skulle aldrig lämna jobbet så . Ni är rädd att något har hänt ? 
Jag kände honom inte , han gick aldrig ur sin roll men han var trevlig . 
Jag vet inte ... Det är konstigt att han inte kom tillbaka . 
- Hamilton ? 
Rappade han ? 
- Du är så rolig ! 
- Var det här det hände ? 
- Lägg av . 
Okej , vad har vi här ? Vi har en gamling som glömmer att ta sina piller och blir förvirrad ? 
- Snackar vi om en virrig gamling ? 
- Nej , det är mer än så . 
Han gick aldrig någonsin ur sin roll . 
Vi har varken namn eller ålder . 
Poliser söker igenom området och tar vittnesmål från gruppen men han verkar bara ha försvunnit . 
- Inspektör Grant . - Ja ? 
Inspektör Sherman . 
Jag är Helen , er nya kriminaltekniker . - En bevistekniker ? 
Är det Nikki ... 
- Braun . 
Så bra och passande . 
En är vit och en är svart . - Minsann . 
- Det var inte min mening . 
Guidningsföretaget gav knappt någonting . 
De hade ett avstängt telefonnummer och en postboxadress . 
Vi måste kolla lokala sjukhus och akutmottagningar . 
Namnet på vår Ben Franklin är Richard Saunders . 
Ni kommer inte att hitta något . Okej . En av mina tidigare existenser hade ett fysiskt tillfredsställande förhållande med mannen i fråga . - Ja , så var det . 
- Det låter coolt . 
Vad menar hon ? 
Hon lekte gömma gurkan med Ben Franklin i ett tidigare liv . 
Vi gjorde mer än delade säng . 
Jag exponerades även för några av hans andra kreativa strävanden däribland skrifter publicerade under pseudonymen " Richard Saunders " . 
Som i " Poor Richard ' s Almanack " . Den är inte bekant ? 
Så vår falske Ben Franklin använder samma pseudonym som den riktige ? 
Ibland kallade han något annat " Richard Saunders " . Hajar ni ? 
- Skämtar hon ? - Nej . 
Vi vet inte vem han är , men han är försvunnen och måste hittas . 
En äldre vandringsguide . 
Hur mycket trubbel kan han vara i ? 
Hej . Vi har kollat efter en Richard Saunders på sjukhusen . Låt mig gissa . Du hade rätt , och det gav inget ? Tack ändå . 
Var det något mer ? 
Du verkade bekymrad över Helen , den nya rättsteknikern ? 
Jag ringde några samtal och hon har förflyttats ofta . 
Trots hennes fläckfria integritet ? 
Vad vet vi om henne ? 
Vetenskap är hennes grej , inte människor . Hennes personlighet har krockat med många överordnade och hon har förflyttats . Mord till sedlighet till kalla fall till oss . 
- Är hon vårt problem nu ? 
- Du vet lika bra som jag att etiketten " svår kvinna " kan ta död på en karriär . 
Hon kanske behöver rätt mentorer . 
- Jag står för det jag sa . - Visst . 
Jag har något här . 
Ben Franklin slängde nyckeln till ett barn . Det kan finnas avtryck på den . 
Be Ethel Merman ta en titt . - Vem ? 
- Bry dig inte om det . 
- Okej ... Hej . - Vad har du hittat ? 
Alla och deras bröder har tagit i den för jag har dussintals ofullständiga avtryck att kolla . 
- Och det gläder dig ? 
- Vi har en svamp bland oss . 
Fläckarna på nyckeln är ett svartmögel , Stachybotrys atra . Det säger inte så mycket för mögel kan växa överallt där det finns vattenskador . 
Men den här nyckeln ... Nycklar består oftast av mässing eller järn men den här är gjord av brons . Ser ni att den är dubbeltandad ? Det är en huvudnyckel , vanlig i byggnader från sent 1700-tal . 
Okej , så vi letar efter en byggnad från kolonialtiden det det finns problem med svartmögel . 
- Jösses . - Vad är det ? 
Ben Franklins möteshus för kväkare . Det byggdes om till internatskola och har varit stängt på grund av mögel . 
- Det verkar vara ett bra gömställe . - Hörni ? 
Skolan brann ner för en timme sedan . 
Jag hämtar Jason och åker dit . 
- Lycka till ! 
- Bra jobbat , Helen . 
- Tack ! Får jag fråga en sak ? - Visst . Har ni hört talas om kryptomnesi ? 
Det är ett fenomen , där folk felaktigt tror att en tanke idé eller upplevelse är ens egen . Ett mentalt tillstånd . 
Antyder du att mina tidigare liv är " ett mentalt tillstånd " ? 
- Det lät illa . - Litegrann . 
Ett tips , de flesta väntar minst en vecka innan de kallar mig galen . 
Jäklar . 
Okej , vi har en accelerator här . Det är definitivt mordbrand . 
Det luktar rena däckfabriken . Vad är det ? 
Latex ? Guiderna bemödar sig verkligen . 
Smink , peruker ... 
- Tjockdräkt ? 
- Japp . 
Vi borde se om den nya tjejen kan hitta några spår . 
Får jag fråga vad du tycker om den nya tjejen ? 
Du ska inte dejta henne , okej ? 
Du fixar inte hennes sjungande . 
Nej . Det är tjejen man kopierade i skolan för att få högsta betyg . 
Hon är väldigt rar . 
Hon gav mig Skittles . 
- Jag fick inga Skittles . 
- Du förtjänar dem inte . 
- Kanske inte . Jag har hittat något . - En bränd madrass ? 
Nej . Se upp nu . 
Får vi låna den ? 
Jag har hittat mycket smuggelgods i madrasser . 
Vi har foton . 
Det var som fan . 
Så nu har vi en mystisk landsfader och en mystisk kvinna ? 
Fotot är inte rent nog för ansiktsigenkänning . 
Inget i databaser eller sociala medier . 
- Och skolan ? 
- Förlåt att ni har fått vänta . Skrivarens färgade bläck tog slut . 
- Är allt det här från brandplatsen ? 
- Jag är noggrann . Ja ! 
Du fick säkert högsta betyg . 
Jag hittade ett fingeravtryck på dräkten . 
Gå till sista sidan . 
Okej . Benjamin Franklins riktiga namn är Owen Maloy . 
Torped för irländska maffian i norra Philly . 
Flera tidigare domar och har varit privatdetektiv men han försvann för tjugo år sedan . 
Det var ett stort maktskifte i maffian då . 
Han kanske tjallade ? Det skulle förklara försvinnandet och den falska identiteten . 
Vem väljer " Ben Franklin " som falskt namn ? 
" Försvinna " och " gömma sig " är helt olika saker . 
Vill du försvinna , lämna delstaten . Varför stanna kvar ? Bilden är tjugo år gammal . Kemi ? Vi har väl fortfarande C:s åldrandeprogram ? 
Jag kör fotot genom det . 
Efterlys honom sedan och kolla upp tjejen . 
Vi måste hitta henne först . 
Maloy har ett uppenbart intresse och en våldsam bakgrund . 
- Händerna på ratten . - Okej , kompis , ta det lugnt . - Vänta nu ... 
Owen ? - Vem mer har du berättat för ? 
- Så det var du i morse ? - Vem mer ? ! 
Ingen . 
Vi trodde att du var död . 
Jag säger inte till någon att jag har sett dig . 
- Jag svär , Owen . 
Jag har en familj ! 
- Ja . 
Kemi . Jag skickade nyss något till dig . 
Det är Charlie McGannon , den nuvarande irländska maffiabossen . 
Polisen och FBI har flera utredningar igång . 
Du sa att det var ett stort maktskifte när vår saknade torped , Owen , gick under jorden . 
Enligt det här blev Charlies far , den gamla bossen , mördad . 
Charlie tog över . 
Inga gripanden gjordes , men Charlie trodde att de egna låg bakom . 
- Tror du att Owen dödade pappan ? 
- Kanske . 
Okej , jag har funderat på den här flickan . 
Om maffian är ute efter killen , varför stanna kvar här ? 
- En enda skulle jag göra det för . - Sidney . 
Flickan på bilderna är Owens dotter . 
Så Owen dödade chefen , försvann och har hållit ett öga på sin dotter . 
- Nu är Charlie efter honom igen . - Killen är en galning . 
Han får Scorsese-filmer att se ut som godnattsagor . 
Vi får larm om att Owen har flytt från en bil i Kensington . 
- Jag hämtar Mike . 
- Fortsätt leta efter Ava . 
Ett vittne såg Owen kliva ur bilen och ett annat såg honom gå söderut . 
- Det är blod . - ... är killen det också . 
- Det där är ett maffiatillhåll . - Och ? 
Någon blir rånad och ringer inte polisen ? 
Han vill inte prata med oss . 
Stället är under övervakning . 
Vi behöver tillstånd för att gå in . 
Tillstånd ? Just det . Vi har ett öppet fall med en saknad maffiatorped . 
Det här är ett känt maffiatillhåll . Vad snackar vi om ? 
Vi kommer att förarga folk utan anledning . 
Nej , vi har en bra anledning . Jag är törstig . 
Kan du slappna av lite ? Ta det lugnt . 
Hur är läget ? 
Kan jag få ett par club soda , tack ? 
- Vi har slut på club soda . 
- Jaså ? 
Är det så uppenbart att vi är snutar ? Va ? 
Det är hans skor , eller hur ? 
Okej . 
Jag försökte , men nu måste vi göra något annat . 
Jag vet inte vad du tänker göra , men gör det inte . 
- Hördu , ta det lugnt ! Allihopa ! Lyssna på mig , okej ? 
Allt är lugnt . 
Jag är polis , från Philadelphiapolisen . 
Såg någon vad som hände med Chryslern utanför ? Med bilen ? 
Någon ? 
Mannen där gnuggar sig i nacken , som om han fått en smäll i skallen . 
Så vad tyckte du om det ? 
" Ingen club soda " ... 
Tjena . Vill du berätta vad som hände ? 
Någon försökte kapa min bil . 
Nej , ingen försökte kapa din bil . 
Din bil står på parkeringen . 
Han heter Owen Maloy , han stack till fots . 
Vi vet att du känner honom . Vi vill veta hur du känner honom . 
Vi tog det tillsammans . 
Är det ni och Charlie McGannon ? 
Ni har känt varandra länge . 
Varför gav han sig på dig ? 
Varför slog Owen dig ? 
Jag trodde att han var död , men i morse visade jag barnbarnen runt och där står han , utklädd till Ben Franklin ! 
Just det . Vad ville han ? 
Killen bredvid Charlie är gamle McGannon . Han var bossen . 
Owen dödade honom och gömde sig . 
Nu vill han veta om någon annan vet att han är kvar i stan . 
Vem mer vet det ? 
Nej ... Owen gjorde ett misstag . Han sa att han har familj . 
Nu vet vi hur vi ska hitta honom . 
Pete , ta det lugnt . 
Ja . Jag har inget mer att säga . 
Kom nu . 
Vi måste hitta Owens dotter innan McGannon och maffian gör det . 
Och de har ett försprång . 
Hur går det med dottern ? 
History Tours skickade allt de hade om Franklin sedan Owen anställdes . Det här är Ben Franklins tidigare rutt . Och det här är rutten som Owen bad att få gå . Ava jobbar nog längs den . 
Vi måste kolla affärsrörelserna . - Hon måste bort från gatan . 
Ms Dufrain ? Kriminalkommissarie Batista . 
Vad händer ? Poliserna sa inget . 
Jag beklagar förvirringen . 
Vi har inte alla bitar på plats ännu . 
Vad kan du berätta om din far ? 
Min far ? Ingenting . Jag har aldrig träffat honom . 
- Han dog när jag var liten . 
- Vi tror att din pappa lever . 
Vi har kollat födelseregistret och upptäckte att din pappa heter Owen Maloy . 
- Du kanske har sett honom så här . 
- Det är Benji . Han är min vän . Han säger åt kunderna att vara snälla mot mig . 
Han är inte min pappa . 
Mamma sa att han blev mördad , för något han inte hade gjort . 
Sa hon vad det var ? 
Ava , vi försöker hitta honom innan något händer honom . 
Håller jag inte öppet , får jag inte betalt . Jag måste gå . 
Jag avråder från det . 
De som letar efter Owen kanske tror att du vet var han är . Men jag kan inte tvinga kvar dig . 
Ring om han tar kontakt . 
- Charlie McGannon . 
- Det var länge sedan . 
- Hur är det ? 
- Mitt kontor . 
- Vad kan jag göra för dig , Charlie ? 
Du har inte förändrats . Jag hörde att du och ditt folk letar efter Owen Maloy . 
- Är det så ? 
- Ja . 
Eller hur ? Det vet du . 
- Hej . 
- Hej . 
Du , det där är Charlie McGannon . 
Du var tvungen att storma in på baren , va ? Nu sitter maffialedaren vid Nikkis skrivbord . Jag ville inte kalla det " stormade " . 
Det där du gjorde är att storma ! 
Nik . Förlåt att jag stör . 
Kan vi snacka lite ? Inte nu . 
Det kan vänta . 
- Är allt bra ? 
- Allt är bra . 
" Nik " ? Doppar du pennan i polisens bläckhorn ? 
- Vad vill du ha av mig , Charlie ? 
- Inget . 
Jag vill att du och ditt folk gör absolut ingenting . 
Owen Maloy är mitt problem . 
Jag tar hand om honom . 
Uppfattat ? 
Vi har känt varandra i många år . Jag har aldrig nånsin jobbat för dig . 
- Se det som en väntjänst . 
- Vi har inte varit vänner heller . 
Lura inte dig själv , Nikki . 
Jag var där . 
Jag behandlade dig som en lillasyster när ditt äktenskap sprack . 
Du ville stiga i graderna och bli chef . 
Och , tja ... 
Du försåg mig med information , men det här är annorlunda . Du bad mig aldrig att titta åt andra hållet då . 
Våra tidigare affärer färgar inte nutiden , Charlie . 
Jag kom hit för att vara artig . Respektfull . 
Ge mig inte anledning att inte vara det . 
Med all respekt , jag är ledsen att du har spillt din tid . 
Vi är poliser och vi ska hitta den saknade personen . 
Okej . Som du vill . 
Vi ses , Nikki . 
- Precis i rättan tid . 
- Det är jag skyldig dig . 
- Vad menar du ? 
Förlåt att jag drog in McGannon . 
Att han hade mage att bara stövla in . Det är inte ditt fel . 
Charlie kom hit på grund av mig . 
- Det finns vissa saker du inte vet . - Vad pratar du om ? 
Jag är en färgad kvinna i ett mansyrke . 
Ingen banade väg för mig , så jag fick göra det själv . 
Charlie var inte lika mäktig då som nu . 
Jag grep honom för droginnehav och fick honom att tjalla . 
- Är han en tjallare ? 
- Han var min informatör . 
Han gav mig information som ledde till många gripanden . 
Charlies gäng har inte lika mycket konkurrens som förr . 
Han satte dit sina rivaler . 
Snabbaste sättet att avsluta ett maffiakrig är att hjälpa en sida . 
Så vad gjorde han här , bad om en tjänst ? 
Maffian är ute efter Owen . 
Enligt ryktet dödade han Charlies pappa och gick under jorden . Du ... Det är okej . 
Vi ska göra vårt jobb och ta Owen levande . 
- Vad är det här ? 
- Intressanta fakta om psykologin bakom tron på tidigare liv . 
Jag har inte bett om din åsikt . 
Det är inte min åsikt . Det är vetenskap . 
Folk har dömt min tro hela mitt liv . 
- Jag klarar mig ändå . Du borde prova . 
- Vad menar du ? 
Har det slagit dig att du förflyttas så ofta för att du anstränger dig för mycket ? 
Fokusera på jobbet . Inte på mig , på jobbet . 
Vi har en försvunnen person med en måltavla på ryggen som behöver oss . 
Förlåt . 
Jag har stängt för dagen . 
Jag är ledsen . 
För vadå ? 
Det är mamma . 
Hon hade samma bild . Hur ... 
Det är vi . 
Det var mitt ex . 
- Är du min pappa ? 
Jag förstår inte . 
Det ... Jag kan inte förklara just nu . 
Det finns inte tid . 
Det finns ett nummer sparat i den . 
Ring om några dagar så kan vi prata när allt har lugnat ner sig . 
Ava ... Att träffa dig var alltid höjdpunkten på min dag . 
Stick härifrån . 
Du måste springa nu ! 
Jag älskar dig . 
Ava är på ditt kontor . Hon vet ingenting . 
Tankarna snurrar . 
Hon träffar sin pappa och sedan blir han bortförd . 
Vittnen sa att han knuffades in i en blå skåpbil . 
Kemi spårade den , men tappade bort den på väg ut ur stan . 
Charlie har honom . Tror han att han sköt hans farsa , så dödar han honom . Inte än . 
Jag fick precis veta att han är här . 
Vem är här ? 
- Se till att han har det han vill ha . 
- Vad har du gjort ? 
Jag gick igenom utredningarna och hittade något att förhöra honom för . 
- Okej , vadå ? - Obetalda parkeringsböter . 
Nikki , det är galet ! 
Hans advokater får ut honom om en timme . 
Missar jag något ? 
Charlies män dödar inte Owen utan hans tillåtelse . 
Hans mobil är bevismaterial . 
Så länge han är här kan han inte ringa och få Owen avrättad . 
Du har rätt . Hans advokat får ut honom om en timme så vi har en timme på oss att hitta Owen Maloy . 
- Jag har redan berättat vad jag vet . 
Jag vet hur svårt det här har varit . 
Som att pappa fick livet åter och sedan dödades igen . 
- Ben Franklin-grejen är så konstig . 
- Inte direkt . 
Om jag var i din fars situation så hade inte jag heller kunnat hålla mig borta från mitt barn . 
Han älskade dig . 
Hamnar han i fängelse om jag hjälper er att hitta honom ? 
Antagligen . 
Men han kommer att vara i livet . 
Han gav mig den här . 
Du gör det rätta . 
Det fanns ett nummer lagrat och jag kunde spåra det . 
De tog I-476 till norr om Allentown innan signalen försvann här . 
- De slog säkert sönder telefonen . 
- De är på väg till Poconos . 
Vänta ... Stugan . 
Vi såg ett foto på en jaktstuga som kan ligga i Poconos . - Ta med Jason och åk dit . 
- Det finns hundratals stugor där . 
Då får vi begränsa sökandet innan de kommer fram . 
- Inte ett knyst från chefen . 
- Du måste lyssna på mig ! 
- Jag dödade inte gamlingen . 
- Kan du få tyst på honom ? 
Vi håller er underrättade . 
Parkförvaltningen och lokalpolisen är redo , men måste veta vart de ska . 
Inga fastigheter står på McGannon eller hans kompanjoner . 
- Om jag bara hade en bild ... - Jag har det . Mike nämnde stugan och jag hittade en kundrecension med en selfie . 
Fotot syns , så jag förstorade det . 
Den digitala kopian finns i din inkorg . 
- Hur kom du på att kolla upp det ? 
- Jag ville hjälpa till . 
Vi har en försvunnen person som är illa ute . 
Okej , vi kollar bilen . 
Ingenting där . 
Det kanske finns ett husnummer ? 
Något där borta ? 
- Herregud ... 
- Begränsar det sökandet ? 
Ja , det gör det . Lite närmare , lite närmare . 
Det är en chinkapin-ek . 
Ser du formen på bladen ? De är avlånga med böljande lober . 
Chinkapin-ek växer nästan bara i och runt Martin ' s Creek . Bra gjort , Helen ! - Meddela Mike . - Okej . - Fan också . - Vad är det ? 
Det är Charlies advokat . 
Owens tid är ute . 
Charlie borde ha ringt nu . 
Jag gillar inte det här . 
Jag beklagar besväret . 
- Lägg av , Nikki . Ge mig min telefon . - Har ingen tagit upp den ? 
- Den är nog kvar hos teknikerna . 
- Jag fick dig dit du är i dag . 
Tro inte att jag inte kan göra det ogjort . 
Jag har din telefon här . Men någon streamade " Masterchef " på den och batteriet dog . 
Tack . 
Ta ut honom . 
Polisen ! 
En nere ! 
Jag har honom på kornet . 
Var är Owen ? 
- Jag ger upp . 
- Owen Maloy ? 
Förlåt . 
Nu ger jag upp . 
Händerna bakom ryggen . 
- Är du okej , Mike ? 
- Ja . 
Irländska maffiastugan . Hur kan jag stå till tjänst ? 
De lade på . 
Jag måste fråga en sak . 
Du kunde ha gömt dig var som helst , gjort vad som helst . 
Varför Ben Franklin ? 
Benjamin Franklin ägde folk . 
Det sista han skrev var ett brev till kongressen om att avskaffa slaveriet . 
Han visade att folk kan förändras och bli ihågkomna för de bra sakerna de gjorde , inte de dåliga . 
Jag gillar den tanken . 
Så det var du hela tiden ? 
Jag kunde inte hålla mig borta . 
Det var din första dag och du gav oss presenter . Du borde få något . 
En kaktus ? 
Butiken bredvid hade inte mycket att välja på . Förlåt . 
Jag är skyldig dig en ursäkt . 
Jag borde inte ha snäst åt dig . Förlåt . Nej , förlåt mig . Särskilt för att du trodde att jag kallade dig galen . 
Jag gillar inte heller att bli målad med den penseln . 
Min mamma är bipolär . 
Det var jobbigt när jag var barn . 
Hennes neurodiversitet fick mig att känna mig galen . 
När jag började i skolan och lärde mig om psykologi och de vetenskapliga orsakerna bakom hennes beteende var det som om ett moln skingrades . 
Allt föll på plats . 
Jag gav dig artiklarna för att visa att jag inte trodde att du var galen . 
Men jag vet att jag måste tona ner det . Nej , nej , jag fattar . 
Vetenskap är din grej . 
Jag följer mitt hjärta . 
Min tro leder mig , men det finns plats för båda . 
Vi har gott om tid att hitta vår väg nu när du är en i teamet . 
En bra första dag . 
Tjena . Du har vänner på mordroteln , eller hur ? Ja , hurså ? Så bra vänner att du kan berätta när rapporten om bilbomben kommer ? 
Du tänker inte släppa det oavsett vad jag säger , va ? 
- Är allt bra ? Vad är det ? - Bara något från tidigare i dag . 
Charlie McGannon . 
Vet du något om deras uppgörelse ? 
Är du arg för att hon känner honom eller för att du inget visste ? 
- Kan jag säga både och ? 
- Ja . 
Nikki kan ta hand om sig själv . Agera inte vit riddare . - " Vit " ? 
Verkligen ? 
- Allt handlar inte om ras . 
Vit riddare är bra . Svart är dåligt . 
Kan en broder rädda dagen ? - Jay ! 
- Ja ? 
Tack . 
Och , allvarligt , släpp det . 
Visst . 
Du är schysst . 
Har du kommit hit för att gotta dig ? 
Jag pratade med Owen om varför han gick under jorden . 
Ryktet sa att han var en förrädare som dödade sin chef , din pappa . 
Men Owen har en annan historia . 
Han säger att han blev kontaktad angående mordet men att han förblev lojal mot farsgubben . 
Din pappa mördades ändå . Owen blev en syndabock medan du stärkte din makt . 
Din egen pappa , Charlie ? 
Det är ett nytt lågvattenmärke . 
Vad tänker du göra med det ogrundade skvallret ? 
Ingenting . Såvida inget händer Ava . 
Eller Owen . 
Kom igen , Nikki . Ta ett glas med mig . Som förr i tiden . 
Kom igen . 
Det här är annorlunda , Charlie . Jag ... Jag ska gifta mig . 
Du har rört om tillräckligt i grytan . 
Gillar fästmannen inte att du har gamla vänner ? 
Han verkade inte vara den kontrollerande typen . 
Mike har inte haft anledning att känna till den delen av mitt liv . 
Det tillhör det förflutna . Nu tror han att jag har hemligheter . 
Har du inte det ? 
- Vi var ett bra team på den tiden . 
- Vi var aldrig ett team . 
Vi hade bara gemensamma intressen under en period . 
Och nu ? 
Nu har vi inte det . 
- Ta hand om dig , Batista . - Det gör jag alltid . 
