Kom igen , rappa på ! 
Bussen väntar inte på någon . 
- Kom igen ! - Kayla , de menar dig . 
Skynda er ! 
Skynda er , ungar ! 
Mamma hade aldrig gjort så . 
Du har rätt , din mamma var smartare än så men till skillnad från henne gillar jag bestraffningar . 
- Kom , vi sätter oss jämte Jordan . 
- Min pappa är så jobbig ! 
- Sitt ner , ungar . 
- Du förtjänar en löneförhöjning . 
Ja , det gör jag . 
Då kör vi . En utflykt till Wagner-institutet . 
Vad gör du , pappa ? 
Okej . 
Okej , då kör vi . 
Jordan , ge den här till Kayla . 
Kayla . Här är ditt vatten . 
Jag behöver inte vatten . 
Sluta hänga runt mig . 
- Lägg ner telefonen och stanna där . - Vad är det ? 
Hallå där ! 
Pappa ! 
Pappa ! 
Varför ? Varför ? 
Hej . Vaknade du precis ? 
Nej , jag har varit uppe i timmar . 
Tränat , tog en smoothie . Toppen . 
Huset börjar se riktigt fint ut . 
- Gillar du det ? 
- Det är jättefint . Jag har bara en fråga . Får han hänga ett basebollträ på väggen ? 
Det användes av J-Roll för att slå en triple mot Cincinnati Reds . 
Hej , Mike . Jag bryr mig inte . 
Mina sportgrejer förvisades till garaget . 
Dina sportgrejer var smutsiga gympaskor och en skateboard . 
- Hej , mamma och pappa . 
- Hej ! - Hej , raring . - Vad gör du ? 
Vaknade du precis ? Min lektion börjar 11.00 och kan ni påminna mig igen varför vi pratar i gryningen ? 
- Mammas idé . 
- Är det mascara ? Har du fortfarande mascara på dig ? Och vems t-shirt är det ? 
Det är inte din t-shirt . 
Jag vet det eftersom du inte går på Penn . 
Vem går på Penn ? Det är Penn State , pappa , och sluta snoka , båda två ! 
Sid , jag älskar dig över allt annat , men du ska veta en sak . Collegekillar är som pirayor . Pirayor vill ha mat . - Collegekillar vill ha ... - Pappa ! 
Jag säger bara , Sid , att du är den bästa tjejen på planeten så alla borde respektera dig , men ... Ölpingis och sånt kan gå lite överstyr , eller hur ? 
Det går överstyr och ... 
Skyll det på ölpingisen . 
Det är rörmokaren . 
Hon är ny . Toppen . Lova bara att ni skyddar er . 
Okej ! Hej då ! 
Älskar dig , Sid . 
Jag älskar dig . 
Jag måste gå . 
- Hollis Braun . - Ja . 
Angenämt . Jag tar över mordroteln , grova brott och försvunna personer . 
Strunta i mustaschen . Jag förlorade ett vad . 
Nej , det är väldigt kommissarie Gordon . 
- Min inre åttaåring tackar dig . - Varsågod . 
Bill har säkert uppdaterat dig . Han höll sig på avstånd . 
Jag hörde det . Avdelningens resultat är verkligen enastående . 
- Tack . - Men Jason Grant-situationen ... 
Ni har ett förflutet , men han är labil . 
Skjuta på parkerade bilar ? Stänga av videon under förhör ? 
Han är Phillys bästa polisman . 
Mitt team fokuserar på att få jobbet gjort . 
Kan du förklara vad ägg har med det att göra ? 
En i mitt team är en shaman . 
En av mina hundar äter sin egen skit om han får , men det får han inte . 
Saken är den att du uppfyller alla mina krav , Nikki . 
- Visst . - Och jag har många . 
Kan du inte kontrollera ditt team , ingen fara , vi löser det . 
Jag är expert på att få problem att försvinna . Förutom den här jäkla mustaschen . 
- Njut av era nya kontor . 
- Tack . 
- Det sa jag inte . - Jösses ! Att du lät honom flytta oss till huvudkontoret . 
Jag hade inget val . 
Han vill hålla ett öga på oss . Särskilt på dig . 
- Okej ... - Oj ! 
Det här får Sidneys studentrum att se städat ut , vilket är bra . 
Det är en fin utsikt . Tror jag . - Vi behöver mycket salvia här . 
- Det är nog inte aktuellt . 
Svara . 
MPU . Mike Sherman . 
- Vänta . Du måste sakta ner . 
- Vad är det ? 
Ja , vi kommer direkt . 
Det var trafikkontoret . 
Läget ? 
De har tittat på alla trafikkameror . Kameran på andra sidan såg bussen köra in , men den kom aldrig ut igen . 
Kom aldrig ut ? 
Bara tio ton buss som försvann ? 
Var David Copperfield här ? 
- Hur många passagerare ? 
- Enligt vår information , 27 . 
Har inte bussarna en GPS ? 
Den är antingen trasig eller avstängd . 
Sätt upp en avspärrning 90 meter på var sida om tunneln . 
Sök igenom alla byggnader . Placera folk på andra sidan också . 
- Mike ? - Ja . 
Vad har du ? Nån har varit här med klätterstövlar . 
Vi borde kolla den kameran . 
- När du säger vi , menar du ... 
- Du . Nej , jag klättrar inte upp där . Jag gör det inte . 
Jag har en dålig rygg . 
I helvete heller . 
Hjälp mig upp . 
- Upp ? - Ja , upp . 
Ursäkta mig ! 
Du , unge man , hjälp inspektören upp här . 
- Ja , sir . 
- Tack . 
- Om jag ramlar dödar Nikki dig . 
- Hon har dödat mig för mindre . 
Mycket imponerande . 
Backa ifall han ramlar , så du inte skadar dig . 
Nån har hackat sändningen . 
Bussen försvann inte . Den kapades . 
Jay , titta där borta ! 
- Hej ! Är du okej ? Prata med mig . 
- Hjälp mig . 
Jag ska hjälpa dig . 
Vad hände ? Min dotter är på bussen . 
Några spår av bussen ? 
Personen som tog buss 447 visste var kamerorna satt . 
Hade de åkt längs 5th Street hade den här sett dem . Hade de kört österut , hade den här sett dem . 
Jag gissar på att de åkte västerut här . 
Allt de behövde göra var att undvika kameror . 
Och försvinna i en stad med 1 300 identiska bussar . 
Men varför skulle nån vilja kidnappa en stadsbuss ? 
Vi vet inte förrän vi vet vilka som är på bussen , förutom barnen . 
När man drar sitt busskort skickar bussen informationen till trafikkontoret . 
Om vi får tillstånd att gå in ... 
- Nej , det tar för lång tid . 
- Vi använder det tunga artilleriet . 
- Hej . 
- Jag har inte tid med det här . 
Inte jag heller . Därför behöver jag dina inloggningsuppgifter . 
Så fan heller . 
Du får ta det med min chef . 
Vet du vad jag hatar mest av allt ? Byråkrati . 
Vi kan sitta här medan jag ringer min chef , som ringer din chef som inte hittar sin chef , för att hon spelar pickleball . Eller så beter vi oss som män och hjälper passagerarna . Du och jag . 
Det finns barn på bussen . 
Tvinga mig inte att skjuta dig . 
Kom igen , kom igen , kom igen . 
Jag är före detta militär . Det var en reflex . 
Om jag hade suttit kvar , så hade jag varit hos henne nu . 
Jag hade gjort samma sak . 
Vi förlorade hennes mamma förra året . I cancer . 
Kayla har gått igenom så mycket , och jag har försökt ... 
Minns du nåt om mannen som kapade bussen ? 
Ja , han bar en mössa . En keps . 
Han är vit , kanske i 40-årsåldern . Det hjälper . Snälla , hjälp mig att hitta mitt barn . Hon har stött bort mig på sistone . Jag borde ha sagt nåt , men jag blev sårad . 
Hon är en toppentjej , kommissarie Batista . 
Det här är hon . 
Okej , unga dam . 
Vad önskade du dig , raring ? 
Att mamma kom tillbaka . 
- Vi ska hitta henne , mr Barosso . - Okej . 
Det är vårt jobb . 
Jag ber om ursäkt . Jason har ett lösenord . 
Jag är inne . 
Så det här är alla barnen . Och det här är alla passagerare som använde ett busskort . 
Kontantbetalningen är nog vår man . 
Ja . Vi har alla passagerares nummer som registrerade sina busskort med ett resekonto . - Alla nummer går till röstbrevlådan . 
- De är avstängda eller blockerade . 
Vi kan inte spåra bussen eller passagerarna . 
Använd AMBER alert . 
Jag har 50 poliser som letar efter en buss . 
Snälla , säg att ni har nåt . 
Baserat på en snabbkoll finns det inga uppenbara kidnappningsmotiv . Inga besöksförbud , inga pågående stämningar . Bara folk som försöker leva sina liv . 
Om det handlar om en lösensumma kommer kidnapparna att höra av sig . 
Jag vill inte vänta . 
Vi har något . Någon såg en av ungarna på Washington Square . 
Åk till Washington Square nu ! 
- Min son var på bussen ! 
- Min dotter är 11 år ! 
Hur tappar man bort en buss ? 
Kommissarie Batista gör allt i sin makt för att få hem era nära och kära . 
Våra poliser tar era kontaktuppgifter . Den bästa hjälpen nu är att åka hem . 
- Nej ! - Du får inte åka hem . Nej . 
Ingen vill gå igenom det här ensam . 
Vi kan väl ordna ett rum ? Eller hur ? 
Jag ska se vad vi kan göra . 
Varsågod . Snälla , en i taget . 
Hej , Baxter . Vilken tur att vi hittade dig på Washington Square . 
Du försökte hitta dina vänner så vad bra att du skippade utflykten . 
Det är bara Wagner-institutet . Jag har redan sett fossilerna fem gånger . 
- Har dina vänner smartmobiler ? 
- Nästan alla . 
Jag frågar det , eftersom vi letar efter kommunikation som kan hjälpa oss att hitta dina vänner . 
- Kommer de att klara sig ? 
- Jag hoppas det . Vi vill identifiera personen som gjorde det här . Men ingen av dina vänner har lagt upp bilder från bussen men du kanske fick ett sms eller ett inlägg ? 
Min son Keith kunde vara riktigt besvärlig . 
Han var smart , men jösses vad han hittade på . 
Jag sa att jag inte blev arg om han gjorde ett misstag utan bara glad om han sa sanningen . Din mamma tycker säkert likadant . 
Enligt pojken som skippade utflykten ska vi kolla " Finstagram " . 
Okej , farmor . Alla säger Finsta , en förkortning av falsk Instagram . 
Många barn skapar de här sidorna med olika namn , så föräldrarna inte ser vad de gör . 
Tror du Sidney har en sån ? 
Jag vet inte , men Kayla Barosso har det . Dottern till mannen som knuffades av bussen . 
Det är @ sexyinpinnk . Pink med två " N " . 
Är hon 12 år ? " Sexig i rosa " ? 
Om vi hittar henne kan du läxa upp henne . 
Ja , hon gjorde inlägg imorse . 
Jag ser bara barn , och ingen av dem är busskaparen . 
Är det en återvändsgränd ? 
Om vi kommer åt live-versionen av fotot kan vi se mer men då måste vi hacka molnet . 
Ingen av mina män är bekväma med det , så nej . 
- Tolv barn , Jay . 
- Jag kanske har ett alternativ . 
- Svart hatt eller vit hatt ? - Gråaktig . 
Briljant . Lite oförutsägbar . Wayne . Hackaren du kände i Afghanistan ? Toppen . Ta in honom . 
Visst . 
Är du galen ? Jag har fredliga avsikter . 
Underbart . Du kan gå på samma sätt . 
Wayne , jag vet att jag svek dig . Jag vet det . Men det är brådskande . 
Som när de läste upp min dom för ett halvår sen . 
Till mitt försvar hade jag problem . 
Du visste om situationen med Keith . 
Nej , efter jag hackade varenda telefon och dator i Afghanistan så svarade du inte ens på mina sms . 
Jag suger . Jag vet . Jag suger . 
Det suger att sitta i ett motellrum med en fotboja som ger mig eksem . 
- Det suger faktiskt . - Ja . 
Jag har ingen mobil , dator eller internet . Jag har bara Cartoon Channel , en ful tavla och ett dött träd . 
Vet du vad det gör med en person ? 
Kom igen , det är inte så illa . 
Du klarade fyra nätter i en grotta med halva talibanerna efter dig . 
Ja , men det fanns en skillnad . 
Jag hade dig . 
Ja . Du drog pappaskämt och gjorde din Eminem-imitation . 
Vilken förresten ... suger . - Nej , 
- Jo . Jag är ledsen att säga det . 
Det är härligt att se dig . 
Och jag kanske kan få ut dig härifrån tillfälligt . 
Skickade våra gamla chefer dig , eller är det din idé ? 
Philadelphiapolisen . Vi har en busslast med försvunna barn , och vi behöver dig . 
- Får jag en dator ? 
Okej . 
Okej . 
Så Jays lilla militärpolare fick ett års husarrest för att ha hackat ryska konsulatet . Hur är det en bra idé ? 
De jobbade för samma säkerhetsföretag . Jay litar på honom . 
- Behöver ni nån som hackar molnet ? 
- Wayne Pascal . Kommissarie Batista . - Exet . 
- Du sa inte att Wayne var en kvinna . 
- Mina föräldrar har humor . 
Hon har också humor , så ni kommer överens bra . 
Vi har ett skrivbord åt dig här borta . 
Jag tar baren . 
Du kan ställa den där borta . Ni hade bra grejer i bevisskåpet . 
Varsågod . 
Stadshuset har fått ett krav på en lösensumma . Vi har fyra timmar på oss att släppa John Maritz som sitter i häktet . 
John Maritz är en idiot . Han hjälper rika att bli av med sina problem . 
Tills han gick för långt . Han fick 16 år för avlyssning och utpressning . 
- Släpps han inte inom fyra timmar börjar de döda passagerare . 
Kommissarie Batista säger att ni är de bästa . 
Bevisa det nu . 
Nej , bussen har inte lokaliserats än , men vi gör allt vi kan . 
Jag vet att min man kommer att försöka spela hjälte . 
Ni är mr Cobis fru , busschauffören ? 
- Snälla , hitta honom . - Varför tog de våra barn ? 
Mina damer och herrar , MPU gör allt vi kan . 
Det här är min Grace . 
Just nu tror vi att era barn är i säkerhet . 
- Hur vet ni det ? 
- Man har begärt en lösensumma . 
- Lösensumma ? 
- Jag har inte råd med det . 
Vänta ! 
Det låter inte som goda nyheter men så länge kidnapparna förhandlar finns det hopp . 
- Vem gjorde det ? - Jag är ledsen . - Att dela detaljer kan äventyra ... 
- Går staden med på deras krav ? 
- Mr Barosso , det är en process . 
- Hon är min dotter ! 
Jag har varit i dina skor . 
Min son , Keith , han blev bortförd . 
Vi fick aldrig tillbaka honom . 
Det är därför som jag jobbar här så ingen annan förälder behöver gå igenom det . 
Så jag hör dig . Det gör jag . 
Jag vet hur du känner , och jag säger inte att det blir lätt . Varje minut känns som ett år , men vi ska få tillbaka era barn ! 
Vartenda ett av dem . 
Lyssna . Du måste ta det lugnt nu när Braun flåsar Nikki i nacken . 
- Lugnt ? " Lugnt " är mitt mellannamn . 
- Sen när ? 
- Säger du att det är mitt fel ? 
- Det är inte motsatsen . Han kommer . 
John Maritz . 
Se så de mäktiga har fallit . 
Det är inte så illa . 
Jag har gått ner några kilo och läser mer . 
Det är avslappnande att slippa folks problem . 
" Folk ? " Det bästa folket hade dig som kortnummer . 
- Jag skvallrar inte . 
- Så ädelt av dig . 
Hur kan vi hjälpa er ? 
Vi undrar om er klient har ett kreativt sätt att lösa sitt fängelseproblem ? 
Jag vet inte vad du pratar om . 
Det skedde en kidnappning idag . 28 personer . 12 av dem är små barn . 
Den försvunna bussen ? Det är ert problem , inte min klients . 
Kidnapparen kräver att han släpps omedelbart så jag säger att det absolut är hans problem . 
John , vi vet att dina konton är frysta men vi tänkte att du har hittat en lösning . Berätta bara , så sticker vi härifrån . Vem betalade du ? 
- Jag betalade ingen . 
- Vem gjorde det ? 
Du är polisen , så du kan väl berätta det . 
Vänta nu , Jason Grant , eller hur ? 
Bara humör , ingen finess . 
Han kunde inte ens få tillbaka sin egen son . 
Jay ! Ta det lugnt ! 
- Vi är nog klara här . - Ja , det är vi . 
Inte illa . 
Vad i helvete lär de ungdomar nuförtiden ? 
- Kom du in på Kaylas konto ? 
- Inte än . Det borde ta cirka 30 sekunder . Hon har ingen tvåstegsverifiering . 
- Ska du hacka hennes lösenord ? - Absolut inte . Få se ... " Första husdjurets namn . " Det här Insta-kontot vet hennes föräldrar om . 
" Saknar min Daisy " , gråtande emoji . Hjärta emoji . " Daisy " . 
Mammas flick ... 
Så , vad gjorde du och Jason i Afghanistan ? 
Det vanliga . Berättade han om när vi kidnappade en kamel ? 
Nej , det gjorde han inte . 
Han utelämnade ett antal saker . 
Jay är som en bok med utrivna blad . Vi står ut med honom för vad vi än missar , så har han världens största hjärta . 
Gamlingar , bingo ! Det måste vara farföräldrarna . 
Kollar metadata , latitud , longitud ... 
Raring ? Vem äger huset på 354 Ardmore Lane ? 
Linda och Mason Hill , och kalla mig inte för raring . 
Inga problem , babe . 
Okej , Hill . Berättade han inte om kamelen ? 
- Nej , det gjorde han inte . 
- Intressant . 
- Inte direkt . 
- En till . 
- Namnet på hennes grundskola . 
Okej . 
Vi är inne . Livebilder . Kör hårt . 
- Och ... där ! 
- Inte nog för att identifiera honom . 
- Toppen . 
- Jag fixar det . 
Snabbt . 
Nej , en strand . 
En skog . 
Nej , en strand . En strand . 
Okej . Nej , vänta . 
Jag är rätt säker på att du är i en park . Hej . 
Ärligt talat , tack . 
Du räddade mig . Det här är ... 
Från vad ? 
Rachel tror att rättsmedicinalverket ger mig ångest så jag försöker meditera . 
Men appen ber mig att hitta mitt lyckliga ställe . 
Är det möjligt att du missar poängen ? 
Nej , poängen är att såvida det inte är akut har jag 15 minuter om dagen . 
Tja ... - Är det kidnapparen från bussen ? - Ja . Du måste identifiera honom . 
Bingo ! Vi har en nödsituation ! 
Kom igen ! 
Varför tog de våra mobiler ? 
Så vi inte kan ringa polisen . Men de vet om det nu . 
Vi måste bara hålla oss lugna . 
Jag vill ha min pappa . 
Jag vet inte ens om han lever . 
- Tänk inte ens tanken , Kay . 
- Han knuffade honom av bussen ! 
Jag är fast med ungarna . Vad händer ? 
Snälla , släpp oss ! 
Håll käften , unge ! 
Okej , vi är på väg . 
Kör förbi stoppskylten ! 
Nästa gång är det din tur . 
C jobbar på en fantombild . 
Philadelphias trafikkontor säger att de inte kan stoppa alla bussar . 
Jag försökte . 
Jag försökte verkligen . 
Är du okej ? 
Om Maritz inte släpps måste jag säga till föräldrarna att om tre timmar kan ett barn dö . Dessutom har Braun läst din akt i detalj . 
Vill du att jag faller vid svärdet ? Nej , vi gör vår grej . 
Det är därför vi är bra . 
Han är smart nog att inse det . Varför är hon kvar ? 
Jag la en hörlur i portföljen som tillhörde Maritz advokat . - Hon spårar den . 
- Varför ? 
Jag tror inte att Maritz gjorde det från fängelset och jag misstänker att hans advokat har kontakt med den som gjorde det . 
- Hur hjälper en hörlur ? 
- Du vill nog inte veta det . 
Det är nåt mer som du inte berättar . 
Kom igen , Nik . 
Varför nämnde du aldrig att Wayne är en kvinna ? 
Inte för att det angår mig längre , men ... 
När du ringde mig och sa att Keith var försvunnen var jag 1 300 mil från alla som betydde nåt för mig . Och jag blev som galen , Nik . 
Jag kunde inte prata eller röra mig . Jag var som paralyserad . 
Wayne sa att hon inte ville att jag skulle resa hem ensam så hon flög hela vägen till Philly med mig , 18 timmar och sen flög hon tillbaka till Bagram . 
Jag vet inte varför jag inte sa nåt . 
Jag visste inte hur du skulle reagera . 
Men jag är skyldig henne en stor tjänst . 
Vart för han oss ? 
Vi försöker , men om han inte släpps har jag en buss med ungar som ... 
- Ja , håll mig underrättad . 
- Vad är det ? 
Chefen säger att staden inte vill släppa Maritz . 
Då har vi drygt två timmar på oss att hitta barnen . 
Min inre röst säger att vi löser det här som alltid men jag vet inte , det här känns annorlunda . Vi fixar det här , okej ? 
Jag har identifierat honom . 
Baz Marsh ! Dömd för mord på en kvinna i Fairhill för två år sen . 
Domen överklagades . 
Han är tidigare dömd för grov vandalism , grov stöld . Oöverlagda brott . 
Det kräket är inte kapabel att planera en kapning . 
- Ta reda på vem som är det . - Har vi en adress ? 
Ja , i mappen . 
Marsh tog bussen . Hur hamnar en snobb som Maritz i maskopi med ett kräk som honom ? 
Med rätt summa pengar kan man få vad man vill . 
- Wayne spårar advokaten nu . 
- Ja , Wayne . Hon verkar påhittig . 
Japp , hon hackade en drönare med tuggummi och en flip-phone . 
- Är ni två en grej ? 
- Vem frågar , du eller Nik ? 
Jag undrar vad ursäkten blir när Braun listar ut att en dömd hackare sitter på våra datorer . 
En brinnande önskan att rädda 28 människor ? Och vi är bara vänner . 
- Typ . - Ja . Exakt . 
Marshs hus borde ligga här på hörnet . 
- Har du hört om att knacka först ? 
- Gjorde jag inte det ? 
Okej , Marsh , vad har du åt oss ? 
En pipborste . Luktar lösningsmedel . 
Rengjort en pistol nyligen . 
Han verkar inte vara typen som får bruna kuvert . 
Eller nån som betalar 3 852 dollar i depositionsavgift . 
Han verkar ha hyrt en affärslokal . 
Första bokstäverna är " CAL " . Adressen är borta , men postnumret är södra Philly . 
Titta här . 
Han visste att barnen skulle vara på bussen . 
- Den jäveln . - Ja . 
Personen som jobbar med Marsh vill åsamka maximal smärta . 
Säg hej . Hej ! 
Jag är kriminalinspektör Jason Grant och jag är ute efter dig . 
Nu sticker vi härifrån . 
Telefonen vi hittade var en kontantmobil med ett nummer som inte funkade . - De undrar om han är identifierad ? 
- Kemi , vad har du på bussen ? 
- De sa södra Philly , eller hur ? - Ja . Så jag matchade bussrutterna med trafikkamerorna . 
Det finns en avvikelse . 
- Det var för 20 minuter sen . 
- Den finns inte på rutten . 
Industriområde , söder om 18th . Vänta . På kvittot står det " CAL " . 
Den gamla Calloway-fabriken ! 
Calloway . Precis här . 
Det tar 15 minuter innan vi är framme . 
Vi har 42 minuter till deadline . 
Vi kan vänta på insatsstyrkan , eller har din bil en dragkrok ? 
Nej , det har jag inte . Hurså ? Strunt samma . 
Jag har en bättre idé . 
Jag tar höger . 
Fan också ! 
Mobilen hemma hos Marsh ? 
Han blev ett problem efter vårt besök . 
Om det här är kidnapparen , vem fan har då passagerarna ? 
Snälla , de är barn . 
Sitt ner ! 
Är det nån mer som har nåt att klaga på ? 
- Hörru ! Chauffören . Upp med dig ! - Nej , varför jag ? - Upp ! Upp med dig ! - Nej , snälla ! 
Sätt fart ! Sluta söla ! 
- Jag har en fru . - Håll käften ! 
Rappa på ! 
Snälla , herrn . 
- Hämta Nik . 
Hallå ! Har ni hittat nåt ? 
Titta , Jay ! 
- Åh , nej . 
- Prata med mig . Ja , de kom igenom här . 
Nik , järnvägen är några hundra meter bort . 
De jävlarna vill hålla dem i rörelse . 
Vi ligger ett steg efter . Barnen betalar priset . 
Det står 31 godståg på bangården . 
- Stäng ner rubbet . 
- Jason , det är omöjligt . Ett tåg avgår var fjärde minut annars stängs hela transportsystemet ner . 
Att söka igenom alla vagnar tar flera timmar . - Ett ögonblick . - Vart ska du ? Vad har du ? 
Maritz advokat är på ett kafé nära hans advokatbyrå . 
Använder han deras wi-fi kan jag hacka hans enheter . 
Nej , allt du hittar godkänns inte som bevis . 
- Det här var din plan . 
- Jag vet det . Jag vill bara inte att det går snett . 
Är du mer orolig för ditt ex , eller att vi inte hinner stoppa kräket ? 
Gör det bara . Okej ? 
- Vad är det för min ? 
- Det här . 
Staden har inte släppt John Maritz inom den angivna tiden . Låt det inte hända igen . 
- Den jäveln . - Ja . 
30 minuter , annars står hon på tur . - Den jäveln ! - Ja . 
Vänta . Ser det ut som insidan av en tågcontainer ? 
- Ja , det gör det . - Ge mig drönarbilder på gården . 
Sätt alla män vi har att söka igenom vagnarna nu ! 
Jag pratade med borgmästaren . 
Mellan den döde busschauffören och att ett barn står på tur , går han med på att släppa Maritz . 
- Gudskelov ! - Tack vare dig . 
Vi gick förbi konferensrummet där familjerna väntar . 
Tack , Braun . 
Vilket för mig till delen som du inte kommer att tacka mig för . 
- Jag vill att MPU drar sig tillbaka . - Vad ? 
Nej ! 
Du ska vara med när frigivningsvillkoren bestäms . Och man retar inte en björn som har ett barn i munnen . 
Jag är glad över borgmästarens beslut men jag litar inte på dem som ligger bakom det här . 
Missade du delen där jag ger order ? 
Du vet att jag har rätt . 
Tolv barn . 
Sabba inte det här . 
Jason och Mike letar fortfarande , men det är en nål i en höstack . 
- Nåt nytt om drönaren ? - Inget än . Men vi kan ha något annat . 
Titta inte på passagerarna , fokusera på kedjan . 
- Kan du zooma in ? - Javisst . 
Den rör sig varannan sekund . 
Är tåget i rörelse ? 
Nej , vagnen står stilla . Bara kedjan rör sig . 
Det står jämte ett tåg som kör förbi . 
Vi räknade hur många gånger kedjan rörde sig , och det var 42 . 
Ett godståg med 42 vagnar körde förbi det . 
Enligt systemet stämmer det in på tåget som körde förbi på spår sju . 
- Ta fram drönarbilden igen . 
- Det är spår sju . 
- Där . På det där flaket . 
- Ge mig ett containernummer . 
- Uppfattat . 
Spärra av den vägen . Vänta på mitt samtal . 
- Jay , var är du ? - Södra sidan av spåret . 
Östra sidan , vid spår sju . Container nummer 7-O-9-1 . 
- Kom hit nu ! 
- Kommer ! 
John Maritz är på väg . 
- Jag har typ fullt upp . 
- Jag hackade advokatens mobil . 
Han representerade vår döde busskapare . 
Jag måste verkligen gå . 
Jag har inte tid just nu , Wayne . 
Och han ringde flera samtal till en klient som också är kriminell . 
Om det är snubben som sköt Marsh så är det samma man som har barnen . 
Vad sjutton är det för oväsen ? 
Bara jag som nästan blev dödad . 
Jag måste gå nu . 
Vänta på mig ! 
Jag går upp . 
- Var är din bil ? Vi måste ringa nu . 
- Precis utanför . 
Nej ! 
Hallå ! 
- Jag har pistolen ! 
- Upp med dig ! 
Händerna bakom ryggen . 
Goda nyheter . Du får sitta resten av livet i en cell med din advokat . Dra åt helvete ! 
- Titta till barnen . - Mår ni bra ? 
Kom igen ! 
- Vi är okej . Låt dem gå . - Inspektör Jason Grant . 
- Spelet är över . Skaffa en advokat . 
- Vi är körda . Kör härifrån ! 
- Nu ! - Maritz ! 
- Där är din pappa . 
Gå ! 
Jag lovade mamma att skydda dig . 
Jag är så ledsen , Kayla . 
Jag lovar att aldrig åka på en skolresa utan dig igen . 
Det gör du säkert . Det är okej . 
Jag älskar dig . Så mycket ! 
- Gillar du football , Nikki ? 
- Det är Philly . Har jag nåt val ? En individ kan göra skillnad , men ett lag kan skapa ett mirakel . 
" Flyg , örnar , flyg ! " 
- Nu avslutar vi det här . 
- Ska bli , chefen . 
Jag kan nu rapportera att kapningen av buss 447 planerades av en advokat som representerar John Maritz . 
Borgmästaren och jag , samt Missing Persons Unit sörjer föraren av buss 447 , Elliot Cobi vars hjältedåd inte kommer att glömmas . 
Angående explosionen som dödade Maritz och hans advokat kommer mordroteln inte att sluta leta förrän vi hittar personen eller personerna som är ansvariga . 
Det var kul så länge det varade . 
Vill du ha en sängfösare ? 
Jag har en fin vintage Gatorade och det finns en ismaskin om du vill ha den kall . 
Jaså ? 
Jag vet inte om jag är redo för Gatorade . 
Okej , då . Du vet var jag finns när du är det . 
Ja ... 
Då så . 
Gudskelov ! 
Maritz begravde många hemligheter för flera mäktiga personer . 
- Nån blev rädd att han skulle tjalla . 
- Det får vi nog aldrig veta . 
Mordroteln ska utreda bilbomben . 
Oavsett , så får barnen sova i sina egna sängar i natt . 
- Vill du göra mig den äran ? 
- Nej . Det brukar vara din grej . 
Se det som en tidig bröllopspresent . 
Du har rätt . 
Det känns bra ! 
Vet du vad som skulle kännas ännu bättre ? En skön ryggmassage . 
- Ett glas vin , ett varmt bad . - Det låter härligt . 
- Säg att det kommer att bli bra här . 
