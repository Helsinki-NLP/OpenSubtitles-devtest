Vi ägnar så mycket tid åt att dölja vilka vi är och att se till att ingen ser vårt rätta jag . Därför är det svårt att minnas en tid då vi gladdes åt att få visa världen vårt sanna jag . 
Imponerande . 
Uniformen klär dig . 
Ser det rätt ut ? Jag fick inte till axelskydden . 
Så där . Perfekt . 
- Vad är det ? - Inget . 
Berätta . 
- Handskarna är felknutna . Ingen ser det . 
- Va ? Fixa det , då ! 
Jag minns mitt första krigsrådsmöte . De var inte lika stora då . Mer privata . - Men Ozai verkar gilla att ha publik . 
- Far säger sig välkomna olika åsikter . 
Jag avråder dig från att prova det . Börja med att observera och lära . 
Så där . 
Hur ser jag ut ? 
Som en prins . 
Varför är vi ur kurs ? Vem bestämde det ? 
- Löjtnant Jee , jag ställde en fråga . 
- Vi fick nya order . 
- Av vem då ? - Av mig . 
Katt och råtta-leken har varat länge nog . Det är dags för en ny strategi . 
Det är jag som jagar avataren . 
Jag leder uppdraget . 
Och jag är amiral . 
Eldfurste Ozai gav mig ansvaret för alla insatser som rör avatarens tillfångatagande . 
Jag välkomnar givetvis din hjälp . 
Jag förväntar mig den . 
Jag behöver alla resurser till hands , oavsett hur små de är . 
Jag tittar förbi sen för att diskutera personalförändringarna som jag vill göra . 
Vad har hänt ? 
Löjtnant Jee , byt kurs igen . 
Hörde du vad jag sa ? 
Byt kurs ! 
Vet du vad straffet för myteri är ? Ja . 
Därför kan jag inte göra som du säger . 
Tänker ni låta det ryggradslösa kräket bestämma över oss ? 
Vi kan inte låta honom ta över efter allt som hänt ! 
De senaste tre åren har vi bara haft varann . Så är det fortfarande . 
Bara vi ombord vet hur det har varit . Zhao förtjänar inte er lojalitet . - Zuko gör det . - Lojalitet ? Med all respekt , general ... Din brorson vet ingenting om lojalitet . 
Annars hade han visat oss , som följt honom dag och natt i tre år , mycket mer respekt . 
Istället får vi stå ut med hans förolämpningar och utbrott . 
Jag vet att Zuko är opolerad . Men du måste förstå att han har varit med om mycket . 
Han vet mycket mer om uppoffringar än du tror . 
Hej , stormästare . Vad bra att ni är här . 
Jag heter Aang och jag vill besöka avatar Rokus tempel . 
Ni förstår , jag är avataren . 
Vi vet det . 
Vänta ! 
Ni ska vara fredens män ! 
Efter honom ! 
Jag är en vän . 
Den här leder till templet . Skynda dig . 
- Han måste vara i närheten ! 
Såja . Lugn , flickan min . 
Fick du vittring ? 
Okej , Nyla . Sätt fart . 
Jag heter Shyu . 
Tyvärr tror stormästaren och de andra att eldfursten är deras sanna andliga ledare . 
De har kommit in på fel spår . 
Tillhörde allt det här Roku ? 
Det är reliker efter tidigare avatarer . Min farfar har bevarat dem . 
Jag måste tala med avatar Roku . Bara han kan hjälpa mig att rädda mina vänner . 
Jag håller dem stången så länge jag kan . 
Kliv åt sidan . 
Stormästare , pojken är avataren . Han utgör världens hopp . 
Kom ihåg avatar Rokus lära . Eld ska inte dominera de andra elementen . Balans ska råda mellan dem . 
Den enda som kan ge oss det är eldfurste Ozai . 
Det är han som ska ena världen , inte avataren . 
Och du anar inte hur mäktig han är på väg att bli . 
För sista gången : Kliv åt sidan . 
Det kan jag inte . 
Då ska du brinna med alla andra icke-troende . 
Vem vågar störa avatarens frid ? 
Det är jag . Aang . 
Brukar man inte buga inför de som är äldre ? 
Och vänta bort blicken ? 
Och hoppa på ett ben ? 
Förlåt ! Jag kunde inte låta bli . 
Det är roligt att se dig , men varför dröjde det så ? Jag trodde att du skulle komma tidigare . 
Avatar Kyoshi sa att jag måste reda ut saker själv . - Att det är en del av resan . 
- Det låter likt henne . 
Kyoshi har alltid varit lite ... Är ni inte alla sådana ? Avatarer är väl inkarnationer av varann ? 
Vi delar samma gnista , men är enskilda individer . 
Jag är olik Kyoshi , precis som du är olik oss båda . 
Vad sa Kyoshi om avatarens roll , till exempel ? 
Att jag måste vara en skoningslös krigare . 
Ja , ibland måste avataren ta till våld och hot , men utöver att vara krigare måste avataren även vara diplomat . 
Kan vi lösa världens problem utan att skada nån ? 
Vi kan försöka , men ett misslyckande får konsekvenser . 
Smärtsamma konsekvenser . 
Men precis som Kyoshi är jag här för att hjälpa dig på din resa . 
- Vad du än behöver . - Det gäller Koh . 
Allt utom det . 
- Du förstår inte . 
- Nej , du förstår inte . 
Koh är en rovlysten ande som kan skada dig värre än du kan föreställa dig . 
Fråga avatar Kuruk . 
Jag har inget val , och tiden rinner ut . 
Han har tillfångatagit mina vänner . Om jag inte gör nåt är de förlorade . 
Snälla . Du har besegrat honom förut . 
Nej , inte besegrat . Jag lyckades bara ta nåt ifrån honom . 
Du kanske har kommit för att återlämna det du stal . 
Ett totem som representerar nåt som Koh behöver och inte kan glömma . 
Smycket tillhörde Ansiktenas moder , en forntida ande som skapade ansikten åt allt levande . 
Det är hennes förtjänst att vi fick identiteter , och hon är Kohs mamma . 
Koh vill ha det alla vill ha . En familj . 
Ett totem ? 
Det kan vi förhandla med . 
Tack , Roku . 
Jag hoppas att du kan rädda dina vänner , men för avataren kan vänner vara en belastning . 
Avataren måste göra omöjliga val , och sätta världens behov före sina egna . Där är Kyoshi och jag överens . 
Lita på mig . 
Det kommer att bespara dig och dina närmaste mycket lidande . 
Vad hände med dem ? 
De är paralyserade . 
Allt kommer att bli bra . 
Du är alltså avataren . 
Så mycket ståhej för ingenting . 
Du måste låta mig gå . 
Allvarligt . Du måste göra det . 
Folk räknar med mig . Du vet inte vad som står på spel . 
Jag har hört att du ska rädda världen . 
Men så här är det . Alla behöver inte räddas . En del av oss har koll på läget . 
Vi har våra eldbändare , jordbändare och vad-som-helst-bändare , och alla vill ha nåt . Alla är beredda att slåss för det . 
Om man är smart , lutar man sig tillbaka och låter dammet lägga sig . Sen kan man plocka åt sig av resterna . 
För min del är världen bra som den är . 
Tiden är ute , avataren . 
Du gjorde det . 
Du fångade honom . 
Räkna gärna . 
Jag litar på dig . Vet du varför ? 
För att vi får dig efter oss om nåt saknas ? 
För att du är så söt . 
Var försiktiga . Det är många som jagar honom . 
Ett gäng jägare har sniffat runt . Dem vill man inte bråka med . 
Vi ses , avataren . 
Snälla , låt mig göra det jag måste göra , så kommer jag tillbaka . 
Mina vänner är i fara . Bara jag kan rädda dem . 
Om jag inte återvänder är de borta för alltid . 
Varför lyssnar du inte på mig ? 
Vet du hur det är att ha ansvar för andra ? - Att ha andras liv i sina händer ? 
Låt mig rädda dem , då ! 
Du kan inte ha varit sån här jämt . 
Vad hände med dig ? 
Jordrikets styrkor är samlade längs den södra kusten . 
Vi försökte flankera dem , men de förlänger linjen . 
En kniptångsmanöver , då ? 
Klipporna är i vägen . De kan kringgå alla attacker . 
Vad tycker du ? 
- Jag föreslår ... - Inte du . 
Zuko . 
Vad tycker du ? 
Hornmönstrat anfall . Omsluta flankerna och lämna en flyktväg . 
Hörde du inte generalen ? De skyddas av klippor på ena sidan . 
Tundrastridsvagnar kan ta sig fram . 
De är jordbändare . Våra stridsvagnar skulle begravas under sten . 
General . 
Vi skulle kunna avancera här . När fiendens eldkraft fokuseras dit , kan vi gå till anfall här och här . 
Hur ska de då kunna gå till reträtt ? 
- Det kan de inte . 
- Då förlorar vi dem . 
Du tänker offra dem . 
Det är en del av krig . 
Vilken division föreslår du ? 
Den 41:a . Det är mest nya rekryter . 
Bra . 
Sånt här lär man sig inte i skolböcker . 
Små pojkar borde veta bättre än att leka krig . 
Det är en usel plan . 
Vad sa du ? 
Jag sa att det är en usel plan ! 
Soldater kommer att dö . För vadå ? 
Det är ovärdigt en Eldnationsofficer . 
- Har du mage att ifrågasätta ... 
Det här kan bara lösas på ett sätt . 
Agni Kai . 
Det är nån där ute . 
- Släpp fram oss ! Vet ni vem jag är ? 
- Självklart . 
Lika väl som vi vet att du har trotsat mina order . Du har varit respektlös mot mig och vanhedrat din far . Det borde väl inte förvåna mig efter allt jag har fått höra . 
Vi tar avataren nu . 
Över min döda kropp . 
Frestande . Men ... 
Yuyan-bågskyttar . 
Ozai var vänlig nog att låna ut dem . 
Det sägs att de kan skjuta vingarna av en eldfluga från tusen stegs avstånd . 
Vart ska du ta honom ? 
Borgen i Pohuai för natten . Sen vidare till huvudstaden . 
Han har väntat länge , och jag vill inte göra honom mer besviken än han redan är . 
- Vi tar det östra passet till Pohuai . 
- Prins Zuko . Vi får se upp för bågskyttarna , men de bevakar säkert ... Zuko ! 
Borgen i Pohuai är ointaglig . 
Varför tror du att Zhao sa att han skulle dit ? 
Det är ett självmordsuppdrag . 
Hela arméer har försökt och misslyckats . 
Dessutom ligger Pohuai innanför Eldnationens gräns . 
- Jag bryr mig inte ! 
- Om Ozai får reda på det ... 
- Men avataren ... 
- Han är borta ! 
För tillfället . 
Just nu har Zhao övertaget , men han kommer att begå misstag , och då ska vi slå till . 
Till dess ... Tålamod . 
Se till att få med allt . Eldfursten vill veta allt om tillfångatagandet . 
Det ska framgå att jag gjorde allt för att få tag i avataren . 
Vi borde få med avatarens tankar också . 
Om inte för eldfursten , så för eftervärlden . 
Då så , avataren . Hade du hört talas om mig innan du tillfångatogs ? 
Snälla . Ni måste släppa mig . 
Det är fyra vakter , inte tre , och både händer och fötter är fjättrade . - Det måste bli rätt . - Oskyldiga liv står på spel ! 
Jag kan inte svika alla igen . 
Inte en gång till . 
Om jag var du skulle jag tänka mindre på mitt förflutna och mer på min framtid . 
Det är inte min framtid som oroar mig . 
Jaså ? 
Jag skulle nog oroa mig lite . 
De dödar dig inte . Då återföds du bara . Då måste vi börja leta på nytt , så du kommer att få leva . 
Men inte gott . 
Blås hur mycket luft du vill . Det förändrar inte ditt öde . 
Vad gör du ? Ta inte med det . 
Vi är lojala söner och döttrar till elden , det överlägsna elementet . 
Bara en sak har stått i vår väg och förhindrat en seger . Avataren . Men idag har vi gjort nåt som ingen annan har lyckats med . 
Vi har fångat avataren ! 
Det här är bara första steget . 
Vi kommer att få utkämpa mäktiga bataljer . Men inte ikväll . 
Vi ska hylla Eldnationen och dess storhet ! 
- Har du allt ? 
- Så klart . Vagnen är fullastad med vin . 
Vilken kväll vi ska ha ! 
Hoppas det blir mindre eldspottande än på Ahns födelsedag . 
Ögonbrynen har nyss vuxit ut igen . 
- Det är lugnt . 
Vem är det ? 
Utlös larmet ! 
Vem är du ? 
Spring först , snacka sen . 
Ta med hela mitt tal , men ändra " lojal " till " trofast " . 
Sa du " lojal " eller " trofast " ? 
Avataren har rymt ! 
- Där ! På muren ! 
- Han får inte nå porten ! 
Avataren ! Stoppa honom ! 
Ta den här ! 
Hoppa på ! 
Ingen eldgivning ! 
Jag behöver avataren levande . 
Vad gör du ? 
Öppna porten ! 
- Gör det ! 
Genast ! 
Öppna porten ! 
Kan du skjuta ? 
Skjut honom . 
Döda legosoldaten och fånga avataren ! 
Nu ! 
Var är de ? 
Kolla där borta ! 
Ser du nåt ? 
Jag har en eka i närheten . 
Vi kan inte gå nånstans när alla soldater är där ute . 
Ligg kvar . 
Du är skadad . 
- Jag tänkte hjälpa dig . - Behövs inte . 
Visst . Som du vill . 
- Vad är det ? 
- Inget . 
Får jag fråga en sak ? 
Gethår eller hare ? 
Din kalligrafipensel . Gethår eller hare ? 
Dina tecken är så prydliga . Jag får inte till mina . Munkarna sa att lemurspillning var lättare att tyda . 
Hör på . Jag borde inte ha tagit din anteckningsbok . Förlåt . Den har varit min räddning . Allvarligt . 
Luftnomadmunkarna ... Alla är borta . Jag hade bara dina anteckningar . 
Jag satt uppe och läste på nätterna . 
Du hjälpte mig . 
Jag menar , de hjälpte mig . 
Gethår . Det är styvare , ger mer kontroll . 
Jag tvingades öva varje morgon . 
Jag fick inte stridsträna förrän jag gjort 100 vertikala och 100 horisontella drag . Samma här ! Men det var för andliga studier . 
Oftast när jag skulle meditera sov jag istället . 
Jag åkte alltid fast . Antagligen för att jag snarkade . 
De där ute tillhör Eldnationen . 
- De är på din sida . Varför flyr du ? 
- De är inte på min sida . 
Men det kommer de att vara när jag fångar dig och ... 
Om jag fångar dig får jag åka hem . Då kan jag inta min plats som tronarvinge . 
Är det nåt du vill ? Att bli nästa eldfurste ? 
Ja , självklart . Det är det alla förväntar sig . 
Gyatso . Han var min lärare . 
Han sa att vi inte kan tänka på andras förväntningar . 
Jag vet . Det är inte så lätt . 
Jag är avataren , och det är det alla förväntar sig av mig . 
Det är det enda jag tänker på . 
Du kanske inte måste vara som andra eldbändare . 
Du kan vara bättre än de . 
Du vet att det eldfursten gör är fel . Du behöver inte vara som han . 
Du kan visa medlidande . 
Hur understår du dig ? 
Jag är Eldnationens kronprins . Jag ska vara en förebild för eldbändare . 
Min far är en stor man . 
Medlidande ? 
Medlidande är ett tecken på svaghet . 
Förlåt . Jag ville inte göra dig illa . 
Andra har redan gjort dig illa så det räcker . 
Gör dig redo . 
Far ? 
Men jag skulle duellera general Li . 
Du är här för att du saknar respekt för vår militär . 
- Det stämmer inte . - Jaså ? 
Även när de kommer på usla planer ? 
Mina planer ! Min strategi . Min militär . Det är det du har förolämpat . 
Förlåt mig . Jag menade inget illa . - Res på dig . - Nej ! 
Snälla ! 
Res på dig ! Bror ! 
Låt bli . 
Han är din son . 
Vi får väl se . 
Res på dig och ta kampen , prins Zuko , så att du kan lära dig att visa respekt . 
Var det allt ? 
Ge mig allt du har ! 
Medlidande är ett tecken på svaghet . 
Soldaterna är borta . Du kan ta dig till din båt utan att nån ser dig . 
Det suger att vara född för 100 år sen . 
Jag saknar mina vänner . 
Som Kuzon . 
Han var bäst . Och han var från Eldnationen . 
Om vi hade känt varann då ... Hade vi blivit vänner då ? 
Du kan gå och lägga dig . Vi håller utkik . 
Vi säger till om vi ser nåt . 
Tack , löjtnant , men jag väntar lite till . 
Du har fel , vet du . Om att han inte bryr sig . 
Zuko bryr sig snarare för mycket , särskilt om alla ombord på skeppet . 
Självklart . 
Löjtnant , har du nånsin frågat dig hur du och de andra fick det här uppdraget ? 
Doktorn har gjort en specialsalva åt dig . 
Det passar inte nu . 
- Jag vill tala med min son . - Han är skadad . 
- Han klarar sig . 
- Men han läker aldrig . 
Doktorn sa att du återhämtar dig snabbt . 
Då är din kropp stark . Det är bra . 
Mentalt , däremot , har du fortfarande brister . 
Du höll igen idag . 
Du kanske tror att du gjorde det av respekt , men det var av svaghet . 
Du måste bli kvitt den svagheten . 
Du måste ge upp den för att bli stark . 
Det är det som gör oss till Eldnationen . 
Därför offrar vi 41:a divisionen . 
Ibland kan de svaga bli starkare . 
Ibland måste man bara ge dem en chans . 
Jag har begått ett misstag . 
Jag har skyddat dig , och det har gjort dig vek som din mor . 
Eftersom du inte kan lära dig läxan här på palatset , kanske världen utanför kan bli en bättre lärare . 
Du ska genast fara härifrån och får inte återvända förrän förrän du har besegrat det största kvarstående hotet mot vår nation . 
Du ska hitta , tillfångata och föra hit avataren . 
Du får inte sätta en fot inom våra gränser innan det är gjort . Annars väntar det strängaste straffet ! - Ozai ! 
Så kan du inte göra ! - Det är redan gjort . 
Och eftersom du oroar dig för 41:a divisionen kan du ta dem med dig som din besättning . 
Fyrtio ... Det är ju vi . 
Ni lever tack vare hans uppoffring . 
Jag ser nåt där ute ! 
Det är han ! Släpp ner repen ! 
- Du är skadad . - Jag mår bra . - Nån borde titta till dig . 
- Jag har varit med om värre . 
Jag tänker inte fråga dig var du har varit , men i framtiden får du gärna meddela om du fortfarande är i livet . 
Det är faktiskt några här som bryr sig om såna saker . 
Givakt ! 
Vår prins har återvänt . 
Vad är det här ? 
De saknade dig på musikkvällen . 
Det är otroligt hur långt vi kan gå för att dölja vårt rätta jag . 
Kanske för att vi inte vill visa folk hur mycket de betyder för oss . Det är lustigt , för vi skulle göra allt för dem . 
Vi skulle resa långt riskera våra liv och bekämpa monster . 
Men det är skrämmande att medge att man behöver nån . 
En del skulle se det som en svaghet . En belastning . 
För finns det nån värre smärta än att förlora nån man älskar ? 
Eller ännu värre ... Gyatso ? 
... att upptäcka att den man älskar har övergett en . 
Kan vi prata om det när jag kommer tillbaka ? 
Självklart . 
Vi får mer tid när jag räddat mina vänner . 
Det är väl därför vi känner ett behov av att skydda oss själva . 
Vi tar på oss en mask . 
Det är inte svårt att förstå varför . 
Det svåra är vetskapen att ibland är masken ens rätta jag . 
