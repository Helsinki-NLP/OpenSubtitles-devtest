Vi måste vara klara senast kl. 14.00 , men bra jobbat . 
- Okej . - Ja . 
Nej , hör på . 
Det kvittar vems getterna är . De måste bort från vägen . 
Lugn , sergeant . 
Försök undvika en internationell incident . 
Okej , herrn med mustasch , gå åt det hållet , tack . 
Herrn med ögonlapp går åt andra hållet . 
Vi löser det fredligt . Låt getterna bestämma . 
- Inga tabbar . 
Bobby ! 
Går det bra ? 
- Hans pass har gått ut . - Får jag se ? 
- Hejsan . - Hej . 
- Det är bara tre dagar . 
Låt dem fortsätta , men bara den här gången . - Det ska fixas innan återresan . - Okej . 
- Freddie . 
- Chefen . 
- Är allt bra ? 
- Jag tar det . - Nej . 
- Jag fixar det . Stanna här . - Ja , sir . 
Jaha . Hej . 
God eftermiddag , sir . 
Ahmed . 
Det bådar inte gott . 
Det var ett otäckt fall . 
- Ni kunde ha ringt . - Det gjorde vi . Flera gånger . 
Till slut bestämde er bror , som den äldsta sonen , att jag skulle sändas iväg för att verkligen inskärpa allvaret i situationen . 
Är min far döende , Ahmed ? 
Hans nåds tillstånd är allvarligt . 
Mina instruktioner är att genast ta er till flygplatsen . 
Era överordnade har gett klartecken . 
Okej . 
Då åker vi . 
Sergeant . 
Kan vi göra nåt , sir ? 
Du för befäl , Charlie . 
Tills jag är tillbaka . 
Välkommen hem , sir . 
- Har du saknat mig , mr Lawrence ? 
Hej , Freddy . 
Eddie . 
Edwina , Edouardo , du är här . Kom . Bra gjort , raring . 
Bra gjort . 
Ge mig en ordentlig kram nu . 
Fint att se dig . 
Hur mår han ? 
- Kasst . - Jaså ? 
Hans kokta fläsk är definitivt stekt . 
Doktorn trodde på ikväll eller imorgon . Du , då ? Hur mår du ? 
Jag har faktiskt ingen aning . Jag är helt ... 
- Hur mår mamma ? 
- Ja , henne får vi hålla ett öga på . 
Hon har nog tagit av pappas mediciner . Ögonen är som navkapslar . 
Okej . 
- Nu samlar vi oss . - Okej . 
Vid det laget var han förstås på pickalurven och spritt språngande naken . 
Han hade glömt att han var i överhusets kammare . 
- Hur tusan ... - Hej , Chuckles . 
- Är du okej ? - Ja . 
- Hur mår han ? 
Är han klartänkt ? - Emellanåt . Till och från . 
När han är med är han ... definitivt med . 
Hej , mamma . 
- Tack och lov . - Herregud . 
Nu blir han glad , även om han inte visar det . 
Ska vi gå ut ? Kom . 
Den första hertigen av Halstead var stenhård . 
Han byggde stället själv . 
Varenda sten . Helt ensam . 
- Pappa ... 
- Snodde sten från det gamla klostret . 
Det är Edward . 
Varför vände du oss ryggen , min son ? 
Tycker du att det är modigt att fara iväg och leka tuffing med dina vänner ? Godset får inte delas upp . Är det förstått ? 
Oroa dig inte för det . Försök vila . 
Och ta hand om din bror . 
Han klarar sig inte utan dig . 
Förstår du ? 
Jag förstår . 
Den tredje hertigen , en elak jävel , dödade 15 fransmän före lunch . 
Han förberedde sig för en duell , men sköt sig själv i foten . 
Den dumma jäveln . 
Doktorn ! 
Eddie . 
... välsignad av den allsmäktiga Gud , Fadern , Sonen och den heliga Anden . 
Må ni alltid bära välsignelsen med er . 
Amen . 
Godset har funnits i släkten i över 600 år , och Freddy lär ... rubbet till jul. 
Vi borde göra nåt åt det . 
Om du hade fått det hade du återförvildat björnar i Berkshire . Än sen ? Jag gillar björnar . 
De lämnar inget koldioxidavtryck och var här före oss . 
Ja , och de äter fan upp en . 
Men det kvittar ju . 
Hela godset går till den förstfödda sonen . 
Det är Freddy som är arvingen . 
Vi kanske borde utföra en kupp . 
Där sa du nåt . 
Ursäkta att jag är sen . 
Där är han . 
Ers nåd . 
Alla smala landsortsvägar ... 
Bra . Kämpa på bara . 
- Jag är strax klar . 
- En kopp te ? Är du okej ? 
Jag fastnade bakom en traktor också . 
Topp . Tipp-topp . - Nej , nej . - Då så . 
Är alla redo ? 
Låt oss få det överstökat . 
Då börjar jag . 
Jag , Archibald Horatio Landrover Horniman , den tolfte hertigen av Halstead , som är vid god vigör , tillkännager detta som min sista vilja och mitt testamente . 
Till Geoffrey Seacombe , för lång och trogen tjänst , överlåter jag besittningsrätt livet ut i grindvaktens stuga . 
Till min fru Sabrina , för hennes lojalitet och trohet under våra lyckliga år tillsammans , lämnar jag ett årligt underhåll som den nya hertigen får överlämna efter behag , samt min älskade labrador Luna . 
Till min dotter Charlotte överlåter jag Endurance , med villkoret att hon seglar världen runt med den inom sex månader . 
Bra , Chuckles . 
Hon får även bundna medel till en summa av 1 000 pund i veckan tills hon gifter sig . Med en man . Jisses . 
Vad gäller resten av min egendom , inklusive min titel , huset och ägorna , den stora vinkällaren , konstsamlingen , yoghurtfarmen och mjölkgården , byn Hetheringham , och fastigheten i södra Frankrike , överlåter jag den härmed till min son ... 
Okej Edward Horniman . 
Jag tror att ... Jag tänkte att alla kunde ... 
Ursäkta . Kan du ta om det där ? 
" Överlåter jag till min son Edward Horniman . " 
Ursäkta . Jag beklagar verkligen . Det måste ha blivit ... 
Han är Edward . Jag är Freddy . 
Ibland kallas jag Fredward , så det kan bli lite rörigt . 
Det verkar ha skett ett misstag . 
Det tror jag inte . 
Jag fattar . Du skämtar . Var det här ... Är det ... 
Har du arrangerat ... Det är ett skämt , va ? Ett sjukt skämt . Det ... 
Jag är den äldsta sonen ! 
Jag ska ärva allt ! - Vad ... 
Vad fan är det här ? - Nej . 
- Det är ett misstag . - Sluta ! 
Lugna dig . 
- Börja inte . 
- Det måste vara ett misstag . 
Jag är den förstfödda sonen . 
Det betyder att jag ärver titeln . 
Det är inte bara jag som säger det . Det står i lagen , för fan ! Det är hämtat från Bibeln , från Gamla testamentet . 
Det är Guds vilja . 
Den förstfödda sonen ärver allt . 
Det är för fan ... Det är förstfödorätt . 
- Förstfödslorätt . 
- Det var ju det jag sa ! 
- Har du hört talas om det ? 
- Givetvis . Men testamentet är tydligt . Godset går till Edward , och titeln har en särskild bestämmelse som tillåter att den andra sonen kan ärva ... 
Ursäkta mig , men jag ger blanka fan i om testamentet är tydligt ! Titta här . 
" Successionsrätt : Det förstfödda , äkta , manliga barnet ... " 
Har du skrivit ut det där ? 
Du kan knipa igen , lady Macbeth . Allvarligt . 
" ... ärver föräldrarnas hela egendom . " 
Huset , titeln , allt , för fan ! Allt ska gå till mig ! 
Varför skakar du på huvudet ? Är du en cocktail ? Sluta med det där ! 
- Mötet ajourneras , Ers nåd . - Freddy ... 
Vi packar ihop nu . Vi får återuppta det här senare . 
Det är över . 
Du kan åka hem nu . Tack så jävla mycket , mr Smithers . 
Mr Burns . 
Nej , inte en chans . Aldrig . 
Den var kul ! 
- Jag ber om ursäkt . - Ingen fara . 
Vi kan gå igenom detaljerna nästa vecka när Freddy har lugnat sig . 
- Han tog det illa . 
- Nu kommer han . Absolut inte . Nej , nej ! 
Det här går fan inte för sig ! 
Ta upp det med Gud ! 
Ta upp det med premiärminist ... Ta upp det med det jävla underhuset ! Eller stoppa upp det i röven ! 
Jag vill ha det som är mitt genom Guds jävla försyn ! Okej ? 
Det var en kniv i hjärtat ! 
Jag faller som London Bridge ! 
Jag har blivit knullad i ansiktet ! 
Påsatt som en hund ! 
Et tu , Brute ? 
Hur gjorde du det , Judas ? 
Ni konspirerar som ormar ! 
Hans nåd vill triumfera . 
Jag visste inget . Jag blev lika förvånad som du . 
Men inte riktigt på samma sätt , va ? 
För första gången på 600 år har släkten avvikit från traditionen . 
Du förbigick din egen storebror ! 
Inte så broderligt av dig . 
Tack , Wham Tam . 
Jag sköter det . Jag kommer snart . 
Hur tror du att jag framstår nu ? 
Hur tror du att det känns ? Hur ska det hjälpa mig att betala mina jävla skulder ? 
Skulder ? 
- Vadå för skulder ? 
- Det låter illavarslande . - Tycker du det ? 
Berätta . 
Minns du Pete Forbes Spencer ? Vi gick på Eton ihop . 
Stort hår , liten kuk , svettiga händer . Kallades Klibbiga Pete . 
Jag minns Pete , men inte hans kuk . 
Tjänade en hacka på fastigheter . Folk köade för att vara med . 
Min miljon växte till 1,5 på tre månader . Det var helt jävla otroligt . 
Sen : en skyskrapa på Maldiverna . Den första . Först till kvarn . 
En , två , tre , fyra miljoner . Pang . 
Och ? 
Tja , sen ... 
Vadå ? 
Sen vändes allt upp och ner . Orkanen slog till . Planet kraschade . Blixten slog ner . 
Torpeden fick fnatt . Vad ska jag säga ? 
Det var inte mitt fel . Gud blåste mig ! 
Var fick du fyra miljoner pund ifrån , Fredward ? 
Från Tommy Dixon . Okej . 
Och vem är det ? 
Vi träffades på avgiftningen . Kokainlangare från Liverpool . 
Han ville låta mig satsa pengarna . Ville ha en del av kakan . 
Så med andra ord är du skyldig en kokainlangare fyra miljoner pund ? 
Jag är skyldig en gangsterfamilj ... 
Du ska nog få , Freddy . 
... åtta miljoner pund . 
Vänta nu . Hur blev fyra åtta ? 
Jag vet inte . Samlad gangsterränta . 
Spelar roll . 
De är gangstrar ! De gör upp reglerna allt eftersom ! 
Allt bra ? 
Tjugofem procent i veckan tills skulden är betald . 
Och de skyr inga medel om man inte betalar i tid . 
Om jag inte betalar den här veckan hugger de av mig kuken . 
Man dör av det . Jag har kollat . 
Jag kan inte ge dig åtta miljoner . 
Du stal min titel , mina pengar och min enda chans att ta mig ur hålet som Gud har grävt åt mig ! 
Och icke att förglömma : Du är skyldig mig ditt liv . 
När du var tre drog jag upp dig ur ankdammen . 
Nej , men jag minns att du ofta tar upp det . 
Jag räddade ditt liv . Nu håller jag på att drunkna , så du måste dra upp mig . 
Freddy ... Jag bad inte om det här . 
Titeln har inget praktiskt värde . 
Verksamheten är olönsam . Det är hål i taket . Staten är girig . 
Lönelistan är hemsk , personalen vämjelig , och du är ett kokainsniffande as . 
Men eftersom du blivit förbisedd och åkt dit med byxorna nere ska jag kolla på det . 
Pappa , vad har du pysslat med ? 
Edward Horniman söker Ahmed Iqbal . Tack . 
Vad kan jag göra för er ? 
Jag behöver en stor summa kontanter den här veckan . 
Hur mycket då ? 
Åtta miljoner pund . 
Kära nån . Herregud . 
Sex miljoner pund . 
Arvet gjorde er till en välbärgad man , men det betyder inte att ni är rik . 
Ni har tillgångar , inte kontanter . 
Berätta . Varför saknar pappas konton större transaktioner de senaste fem åren ? 
Vi diskuterade aldrig hans privata utgifter . 
Okej . 
Obligationer och aktier , då ? 
- Det finns inga . - Va ? 
Det kan ha funnits annat som vi inte tog upp , men det vet jag förstås inget om . 
Det lät ganska kryptiskt . 
Ni kan sälja Gainsboroughn , men om ni ska få ut det rätta värdet lär det ta flera månader . 
En advokat i London har gjort en okonventionell trevare . 
Hans klient är intresserad av att köpa Halsteads herrgård . 
När nån dör samlas gamarna . 
Ganska fräckt , va ? 
Vad heter han ? 
Den potentiella köparen vill vara anonym i nuläget . 
Men advokaten uppgav att han är beredd att betala långt över marknadsvärdet . 
Det kan alltså ge en ansenlig summa , men bouppteckningen och kapitalvinsten måste räknas med . 
Hälsa dem att jag är beredd att lyssna om han är aggressiv och snabb . 
Förlåt om jag påtalar det uppenbara , men jag skulle försumma mina plikter om jag inte påpekade att Halstead varit i släktens ägo i flera generationer . 
Sedan 1550 . 
Men som sagt : Jag måste ha pengarna den här veckan . 
- Ordna ett möte , är du snäll . - Uppfattat . 
Ursäkta att jag stör . 
Jag ska presentera mig . 
Jag heter Susie Glass . 
Hur kan jag hjälpa dig ? 
Jag gjorde affärer med din far . 
Ursäkta , men pappa var inte direkt känd för sitt sinne för affärer . 
Jag har vissa intressen som jag måste diskutera med dig . 
Som vadå ? 
Det är enklare att visa dig . 
Jag gillade din far . 
En riktig gentleman . 
Lite excentrisk , men adeln är ju det . 
Det måste ha varit en chock att få ärva allt . Huset , titeln ... 
Värre saker har hänt . 
- Nämnde han intäkterna från gården ? Hade de varit betydande hade jag vetat om dem . 
Det beror väl på vad man ser som " betydande " . 
Han drog in fem miljoner pund per år . Plus vinstutdelning . 
Ursäkta ? Fem miljoner pund ? 
Inte för yoghurt och hamburgare , väl ? 
Följ med mig . 
Vad pågår där nere ? 
Vad i helvete är det som pågår ? 
Den brittiska cannabismarknaden är värd över sex miljarder per år . 
Vi har erövrat en ansenlig del av den , men odlingarna tar plats . Där kom din far in i bilden . 
Mot en generös ersättning lät han oss hållas utan att lägga sig i . 
Det finns få egendomar på 6 000 hektar där man i tysthet kan göra vad man vill . 
- Vad heter den här , Jimmy ? 
- Frisian duck . 
Ganska poppis just nu . 
Det här är Jimmy . Han har varit produktchef här i ... Hur länge är det nu ? 
Tre år . Så länge har jag bott under ditt tak . 
Kul att äntligen träffas ! 
Du tillhör familjen . 
Förutom att du typ är en hertig eller nåt . 
Trevligt att äntligen träffas . 
Jag antar att pappa fick ungefär tio procent per år . Det vore inte mer än rätt . Då måste ni dra in 50 miljoner per år . 
I runda slängar . 
Och du sa att ni har en ansenlig del av marknaden . Jag antar att det betyder hälften eller mer . Då måste det här vara en liten kugge i ett större maskineri . 
Ni måste ha dussintals såna här ställen . 
Din pappa brydde sig aldrig om verksamhetens upplägg . 
Jag är nyfiken av mig . 
Det räcker att du vet att vi har ett avtal , och att du som ny hyresvärd får en stor summa pengar varje år i utbyte mot att låta oss hållas . 
Problemet är att jag kanske måste sälja huset . 
Vi föredrar nuvarande upplägg . 
Jag beklagar om du hamnar i kläm , ms Glass , men jag kanske inte har nåt val . 
Jag förstår , Ers nåd . 
Vad händer om jag vill omförhandla ? 
Om du menade allvar med att sälja godset blir det en utmaning för oss . 
- Juridiskt sett kan ni inget göra . - Nej . 
Juridiskt sett kan vi inget göra . 
Var det ett förtäckt hot ? 
Absolut inte . 
Det är mycket att smälta . Jag förstår det . 
Vanligtvis brukar man diskutera sånt här på förhand . 
Och vanligtvis tar den viljesvaga , arbetsskygga arvingen emot pengarna och fogar sig som en duktig liten pojke . 
Så skulle jag inte uttrycka det . Men ja . 
Låt tanken ligga till sig . Vill du ha skjuts tillbaka ? 
Nej , tack . Jag går . 
Ers nåd . 
Hej , Geoff . 
Jag hittade henne vid sjön . Tänkte ta henne till huset . 
Jag vill gärna prata med dig om du har tid . 
Jag brukar ta en kopp te så här dags . 
Perfekt . 
Hur länge har du jobbat här ? Är det 20 år nu ? 
Jag är inte bra på årtal , men ni och er bror var små . 
Du har varit otroligt lojal mot pappa . 
Han gav en bråkstake en chans . 
Det behövde han inte göra , men det gjorde han . 
Jag vet att inget händer här utan att du vet om det . 
Det kan man säga . 
Så jag antar att du har viss koll på läget . 
Det kan man också säga . 
- Mjölk och socker ? - Tack . 
Ni har visst träffat ms Glass . 
Så jag gissar att även ni har koll på läget . 
Hur inblandad är du ? 
Jag ser till att hålla mig utanför . 
Sex tusen hektar håller mig sysselsatt . 
Särskilt när du tar hand om alla skadade djur du ser . 
Det är som ett zoo . 
Charlie blev påkörd av en bil . Sarah-Jane flög in i ett fönster . 
Och den här lilla krabaten har brutit benet . 
Är det en räv ? 
Ska du inte gallra ut rävar ? 
Var det nåt särskilt ni ville fråga ? Ja . 
Pappa var nöjd med läget , men jag är inte lika bekväm med det . 
Det kan bli svårt . 
De är inga skojare , ska ni veta . 
Borde jag ta pengarna och knipa käft ? 
Det funkade för er far . 
Nu har de rotat sig . 
Saken är att jag sitter i en knivig sits . Och av olika anledningar behöver jag deras hjälp . 
Det kan de ge er . Men det kostar . 
- Vad vet du om dem ? 
- De är farliga jävlar . 
I grunden är de affärsmän . 
Så länge de tjänar på det är de beredda att lyssna . 
Var försiktig . 
De ser rumsrena ut , men låt er inte luras av fasaden . 
Hej , Ahmed . Edward Horniman . 
Jag ska inte sälja huset . 
- Tack , Bradley . 
God morgon , Chuckles . Edwina . 
- En kopp te ? 
- Hinner inte . Jag ska med tåget . 
- Är du klädd för jordenruntresan ? - Ser det så ut ? Nej . 
Mamma övertalade mig att avsluta studieåret . 
Det låter vettigt . 
Det är Freddy hon ska oroa sig för . 
Oroa dig inte för Freddy . 
Honom tar jag hand om . 
Behöver du bärhjälp ? Av dig ? Herrn i huset ? 
Bradley . 
Javisst , Ers nåd . 
Lycka till , Chuckles . 
Ers nåd . 
Sätt fart , Bradley . 
Jacky ! Kom hit . 
Det är hertigen . 
- Hejsan . 
- Jag måste snabbt få in åtta miljoner . 
Det var en stor siffra . 
Min bror har skulder till en langare i Liverpool . 
- Har du ett namn ? 
- Tommy Dixon . 
Jag vet vem det är . 
- Hur mycket är ränta ? 
- Hälften . 
Det var hårt . 
Räntan framgick inte när min bror tog lånet . 
Och mina möjligheter att få ihop det som krävs är starkt begränsade , med tanke på vårt avtal . 
Jag ska se vad jag kan göra . 
Hur mycket kan du få ihop ? 
Vet inte . Jag jobbar på det . 
Om du kan fixa fram fyra ska jag se vad jag kan göra med resten . 
Jag återkommer . 
Vad tror du ? 
Jag vet vem Tommy är . Och hans bror , Gospel . 
Ett par knarklangare som har Gud på sin sida . 
- Stygga ? 
- Ja , men inte utöver det vanliga . 
Du kan klämma åt dem . När de fattar vem pappa är . 
Var finns de ? 
Fiskhallen . Bakom makrillen . Det är deras fasad . 
Kom nu , Jacky ! 
Gå tillbaka du . 
Elmo , inkommande . 
Gör dig inte illa . 
Jag heter Stevens . 
Jag är assistent åt privatpersonen som vill köpa Halsteads herrgård . 
Jag måste säga att min klient blev besviken när er advokat sa att ni dragit er ur förhandlingarna innan han fått chansen att kontra med ett mer attraktivt erbjudande . 
Det oaktat undrar min klient om ni kan tänka er ett möte öga mot öga . 
Och vem är din klient ? 
Om ni följer med mig kan ni ses redan nu på förmiddagen . 
Tack , men läget har förändrats . Jag ska inte sälja huset . Mr Lawrence . 
Min klient förstår att det här är en olägenhet för er . 
Därför vill han ge er ett erbjudande . 
Tvåhundrafemtio tusen brittiska pund . För er tid . 
Utan återbetalningskrav , så klart . 
Vill ni följa med mig ? 
Fin piggvar . Två och ett halvt kilo . 
Inte illa för en vild fisk . 
Ska du titta eller köpa , vännen ? 
Ingetdera . Jag söker dig . 
Jag heter Susie Glass . 
Bobby Glass vältaliga och eleganta dotter . 
Jag respekterar Bobby . 
Det gör alla . 
Kan vi talas vid ? Angående Freddy Horniman . 
Tjugofem procent i veckan . Tills skulden är betald . 
Vi går upp . 
Din pappa har tydligen åkt på en förkylning . 
Hur länge har han kvar ? 
- Han har suttit av fyra år av tio . 
Jag har bara hört bra saker om dig . 
Jag trodde inte att braja var värt besväret . 
Skrymmande , små vinster ... 
Men du verkar ha koll på läget . 
Vi har aldrig sysslat med koks , så vi konkurrerar inte . 
Jag förstår inte vad du har för koppling till den där sprätten . 
Jag har affärsintressen som kan äventyras av hans lilla skuld . 
Jag ville höra om det gick att lösa . 
- Åtta miljoner är mycket pengar . 
- Men 100 % av inget är inte ett skit . 
Vi vet båda att du inte får hela summan , så var lite realistisk . 
Vad händer om jag får fram de ursprungliga fyra till slutet av veckan ? 
Jag kan inte skriva av fyra miljoner i ränta . 
Kan vi inte se det som en investering i din verksamhet ? 
Nej , jag söker inte investerare . 
Men jag försöker hitta ett sätt att lösa det här på nåt sätt . 
När får jag de fyra miljonerna ? 
Du kan hämta dem på fredag , och få White Widow för en mille på köpet . 
Okej . 
På ett villkor . 
Han måste be om ursäkt . Och erkänna att han är ett kukhuvud . 
Uppfattat . 
Jag vill spela in det för eftervärlden . 
Det ska efterlikna en video jag har . 
Okej . 
Det finns många sorters videor . 
Det är inget otäckt . 
Då så . Om du får fyra mille och brajan och videon med en ursäkt ... Är det lugnt sen ? 
Ja . Fixar du allt det så är det kolugnt . 
Tack , Jeffrey . 
Sir , hertigen av Halstead , Edward Horniman . 
God morgon . 
Ett nöje , Ers nåd . 
Stanley Johnston . Med ett " T " . 
Du undrar säkert varför jag så gärna vill köpa ditt familjegods . 
Ja , faktiskt . 
Tack , Stevens . 
Sanningen är att det är ett praktexempel på William Kents arkitektoniska filosofi . Han var en tusenkonstnär . Och mästerlig . 
Är du bekant med hans filosofi ? 
Handlade den inte om försoning mellan det vilda och det förfinade ? 
Ett värdigt intresse som vi delar . 
Människor kan överleva i djungeln eller existera i en djurpark . 
Få inser betydelsen av den paradoxala försoningen mellan alternativen . 
Det krävs en sällsynt individ som förstår hur listig och aggressiv man måste vara för att förvärva en egendom som din . 
Ditt hus är ett bevis på den här kulturens syntes . 
Förfining med aggression . 
Den första hertigen förstod den principen , precis som jag . 
Därför ska jag erbjuda dig en obscen summa pengar för ditt lantgods . 
Det låter övertygande . 
Men det kan lika gärna övertyga mig att inte sälja . 
Ska vi spela eller prata ? 
Dricker du vin ? 
Värde härstammar från det som nån är beredd att betala för nåt . 
Om jag säger att det är värt så mycket , så är det så . För mig . 
Det var en rejäl siffra . 
Och jag uppskattar dina ansträngningar . 
Men jag har ändrat mig . Godset är inte till salu . 
Tack . 
Jag hoppas att du inte misstycker till mitt sätt att dricka vin . Jag går emot traditionen och häller upp och filtrerar vätskan . Rengör flaskan från avlagringar . Sen hälls vinet tillbaka för att avnjutas ur sin ursprungliga boning . 
På tal om boningar ... Jag är beredd att höja siffran markant . 
Varför inte låta mig befria dig från din arvsbörda ? 
Det kanske förvånar dig , men jag uppskattar den paradoxala välsignelsen och förbannelsen av ditt upplevda privilegium . 
Jag uppskattar det , men tajming betyder allt , och det här är fel tidpunkt . 
Stevens , var så snäll . 
Mr J. 
- Tack . 
- Så gärna . 
Smaskigt . 
Romanée-Conti från 2002 . 
Gillar du DRC ? 
Jag föredrar Bordeaux . 
Men pappa var förtjust i bourgogneviner . 
Han samlade på DRC . 
Har du provat en från - 82 ? 
Det finns tydligen bara sex lådor kvar i hela världen . 
Åtta , faktiskt . 
Två tillhör kronogodset , en tillhör ärkehertigen av Moldavien och resten står i vår källare . 
Liksom två lådor av den från - 45 . 
Frestelsen blir för stor . 
Låt mig åtminstone få köpa vinet . 
Jag lovar att vara generös . 
Vinsamlingen , då ? 
Den kan ge tre , men det kommer att ta tid . 
Det kan jag svårligen skiljas ifrån . 
- Ers nåd . 
- Mr Stevens . 
Nu kör vi . 
- Det är pappas vinsamling . - I pappersform . Perfekt . 
Det och pengarna i kassaskåpet borde täcka Freddys skulder . 
Om samtalet med mr Dixon gick bra . 
Han hade några förbehåll . 
Han godtar fyra , om det är kontant och imorgon . 
Från åtta till fyra . Imponerande . 
Se det som en gest av välvilja . Från min sida . 
Är allt bra ? 
Inte direkt . 
Eddie , Eddie ... 
Edwina , lyssna på mig , okej ? Killen är tvåfaldig världsmästare i tungvikt . 
- Hur mycket har du satsat ? 
- Alltihop . 
Det är bergsäkert . Jag träffade tränaren . 
Vad heter vadhållaren du använde ? Svara . 
Det finns inga vadhållare . Fajten är exklusiv och inofficiell . Det är V-V-VIP . 
Men hur kunde du satsa nåt utan en vadhållare ? 
- Genom en vän till en vän . 
- Vad menar du ? Vem då ? 
Pete . Hans polare satsade fem mille . - Jag fick vara med . 
- För helvete . Klibbiga Pete ? 
- Har du inte lärt dig nånting ? 
- Han vill gottgöra mig . 
Segern är kassaskåpssäker . Det är Joey Bang * Bang . 
Säg att det var ett misstag . Be om ursäkt och ta tillbaka pengarna . 
Jag måste sluta . Det är mobilförbud här . Så exklusivt är det . 
- Lyssna på mig ! 
- Jag lägger på nu . Älskar dig . 
Ikväll blir det fajt . 
Härligt ! 
- Vi måste ta reda på var han är . 
- Jag känner nån . 
- Läget , Suze ? - Jacky . 
Ers höghet . 
Jack . 
- Har du pengarna ? 
- Ja . Här . 
- Två hundra , va ? - Ja . Jag kan inte lova nåt . 
Jag snackar med dörrvakten , så får vi se . 
Vänta här . 
Din bror verkar välfungerande . Måste vara trevligt . 
- Det är han inte jämt . 
- Vad har han för last ? 
- Kuken . 
- Vad gör han med den ? 
Det vanliga . Men mycket av det . 
Jag lyckades fixa två biljetter . 
Men hör på . Fajten sker helt utanför protokollet . 
Resultatet får inte spridas , för båda är världsmästarboxare . 
De kan förlora sin rankning . 
Och Suze , inget bråk . Mitt namn står på spel . 
- Okej . 
- Ha så kul . 
Okej . Nu tar vi tillbaka pengarna . 
Det är inte ofta de ordnar sånt här . 
De där har flugit hit från Vegas . 
Gypsy Kid är populär på andra sidan Atlanten . 
Joey Bang * Bang drar folk . 
Vi har amerikanerna . Och så albanerna och kineserna . 
Och ryssarna , som glatt sitter bredvid ukrainarna . 
Och så resandefolket . 
Ge honom bara ! 
Inget samlar folk som lite blod i ringen . 
Det lär omsättas 50-100 miljoner pund här ikväll . 
Ja . Och några av dem är mina . 
Psykologi , baby . 
Edwina , hur fan kom du in ? - Pengarna . - Va ? Freddys pengar . De är mina . 
Det är för sent . Fajten har börjat . 
- Eddie , jag har läget under kontroll . 
- Dig tar jag itu med sen . 
Leta reda på vadslagaren och ta tillbaka pengarna . 
Slappna av . Bang * Bang kan inte förlora . 
Han gör mos av honom . Du sabbar stämningen . 
Det är fajt ikväll ! 
- Kan vi ta det här sen ? Jag vill titta . 
Du vet inte om det , men du har klivit in i en främmande värld . 
Nån som inte tål att bli besviken ska ha de där pengarna . 
Förlåt , men det lät som ett hot . Det är inte mitt bekymmer . 
Det kommer att bli ditt . 
Din bror satte pengarna på Joey . 
Om han vinner dubblas pengarna . Om han förlorar är pengarna inte hans längre . Det kan ingen göra nåt åt . 
Ta det lugnt . 
Susie Glass vill prata med dig . 
- Det här är inte över . - Visst . Dra åt helvete med dig . 
Tack , Roger . 
- Hur gick det ? 
- Inte så bra som jag hade velat . 
Sätt dig , ta en drink , titta på fajten . Vi löser det . 
Det här fixar du , Bang * Bang ! 
Vadå ? Vad är det ? 
Han är en svindlare . 
Vad menar du ? 
Han satsar aldrig pengarna . 
Han ger sig på snobbarna . Bara de privilegierade . 
Han skyddar sig med plastgangstrar som han beblandat sig med , och din sort vågar inte protestera . 
Du satsade aldrig pengarna . 
Det är en allvarlig anklagelse , Ers nåd . 
Reglerna för vadslagning är ganska enkla . Förlorar man , måste man betala . 
Vad säger du , John ? 
Jag tycker att du ska dra hem till ditt lantgods och runka av din spaniel . 
- Släpp mig . 
- Passa dig , din sprätt . 
Vi vet var du bor och kan hälsa på . 
Du skämmer ut dig . 
Du tillhör inte armén längre . Och du har inga bevis . 
Varför ligger han på golvet ! Lyft upp honom ! 
Nej ! Helvete också ! 
- Några framsteg ? - Nej . 
Vi måste gå . Nu . 
Får jag tala med honom ? 
När det har lugnat ner sig . 
Känner du igen namnet Stanley Johnston ? 
Nej . Hur så ? 
Det var honom jag sålde vinet till . Han vill köpa godset . 
Summan han erbjöd tyder på att han känner till verksamheten . 
Vad hette han ? 
Stanley Johnston . 
Med ett " T " . 
Vad sa du till honom ? 
Att jag inte vill sälja . Bra . Det var rätt svar . 
Titta på det här . 
Vad är det ? 
Texten till en sång Freddy ska sjunga när han överlämnar pengarna . 
Och han måste dansa . Som en höna . 
- Som en höna ? 
- Ja . 
Varför det ? 
För att Tommy Dixon vill ha en ursäkt , förståeligt nog . 
Det är dags . 
" Jag är en sprätt som tabbade sig , lian , lian , lej . 
Att tabba sig har blivit en grej , lian , lian , lej . 
Men en kuk-kuk här och en kuk-kuk där ... " 
Hur gammal är Tommy Dixon ? 
Vi kommer lindrigt undan . 
- Ska vi räkna dem ? Jag har inte kollat . 
- Det är lugnt . 
- Säkert ? 
Det tar bara en stund . 
- Nej , vi drar . 
Okej . 
Han verkar vilja be om ursäkt . 
Vill du ha en ursäkt ? 
Vet inte . Vill jag det ? 
Ja . Så får vi ett avslut . 
Blanket ! 
En Klibbig Pete . 
Jag ville bara be om ursäkt från djupet av mitt hjärta . 
Fint , va ? 
Du fick pengarna och jag har bett om ursäkt . Är det lugnt nu ? 
Jag vet inte . 
Är det lugnt , Edward ? 
Ja . Det är lugnt . 
- Du sa att ni skulle prata med honom . 
- Det gjorde vi . 
Oroa dig inte . Vi gjorde honom en tjänst . 
Vi straffar hunden , inte mannen . 
Vad ska det betyda ? 
Han har en hund i sig som han inte kan styra över . Vi fick göra det åt honom . 
Vet du vad människans stora utmaning är ? Nej . 
Men om jag läser mellan raderna ... För mycket hund , för lite man ? 
För mycket otränad hund . Och vi är hundtränare . 
Helvete också ! Jag har missat tio på raken ! 
Vikten är fel . De flyger för fort . 
Skjut inte på målet den här gången . Skjut en meter framför . 
Det är ju det jag gör . 
Försök att missa framför , då . 
Där satt den ! 
Född till att döda . Bra där . Edwina . 
Ja , tack , mr Lawrence . 
- Wham Tam . 
- Edwina . 
Hur gick det med Pete ? 
- Jag fick tillbaka pengarna . - Va ? Hur då ? 
- Han satsade dem aldrig . 
- Vad menar du ? 
Han satsade inte pengarna . 
Den jävla ... 
Men mr Dixon har gått med på fyra , så allt är klart inför imorgon . 
Det var som fan . Hur lyckades du med det ? 
Fyra miljoner mindre . Herregud . Jag skulle suga av honom för fyra . 
Bra att veta . 
Men det finns en liten hake . 
- Vad menar du ? 
Du ska säga att du är ett kukhuvud . 
Ska jag ... 
Visst . Jag är ett kukhuvud . 
Så . Skitenkelt . Inga problem . 
Vad bra . 
Alla tycker det ändå . Han gör det . Pete gör det . 
Och pappa . Annars hade han inte gjort mig arvlös . 
Tycker du att jag är det ? 
- Du har varit lite av ett kukhuvud . 
Du är inte alltid det . 
Det är ju jävligt ... 
Geoff , är jag ett kukhuvud ? 
Tackar . Wham Tam ? Är jag ett kukhuvud ? 
Alla män är det , Freddy . - Visst . Var det nåt mer ? 
Han vill att du ska dansa och sjunga ursäkten . Så här . 
- Han har en hönsdräkt . 
- Ja . Det också . 
Okej . 
Jag är en höna . Kackel , kackel , förlåt . 
Så där . Mer , då ? 
Han vill filma det . 
Nej . 
Jag vägrar . Aldrig i helvete . 
Nyss var du beredd att suga av honom . 
I enrum , ja . 
Han ska filma det . 
Nej , det ska han fan inte ! 
Jo , det ska han . 
Du bad om min hjälp . Nu får du den . 
Inte för att du räddade mig när jag var tre , utan för att du är min bror och det är sånt bröder gör . 
Därför måste du göra exakt som jag säger hädanefter . 
Om det betyder att du ska dansa som en höna , så gör du det . 
Då dansar du inte som en strippa , en björn eller en jävla ballerina . Du dansar som en höna . 
Är det förstått ? 
Ska du ta återstoden av min värdighet också ? 
Har du förstått , Freddy ? 
Ja , Ers nåd . 
Vilket ställe . 
Thomas . Bakdörren , sa jag . 
Tjänsteingången . Det gäller ju trots allt en tjänst . 
Jag gick ner från åtta till fyra . Nog kan jag använda huvudingången . 
Kom , då . 
Hörru , grabben . Glöm inte dräkten . 
- God dag , herr Dixon . - Tjena . 
Tack för att du kom . Vi vet att du är en upptagen man . 
Det var en fin biltur . 
Vackert landskap . 
Är det till mig ? 
- Som utlovat . Vill du räkna dem ? 
- Nej , det kan Jethro göra . 
Jezza , din tur . 
Hörru ! Grabben ! 
Får han låna skrivbordet ? 
Javisst . Slå dig ner . 
Han har tvångssyndrom . Han är trög i starten , men sen är han ostoppbar . Då så . Ska vi köra igång ? 
Hör på , Tommy . Den här hönsgrejen ... 
Alltså ... Jag kan bära dräkten och dansa , för att visa hur uppriktigt ledsen jag är för det här . Men du får dina pengar , du får ditt roliga och jag får kräla ordentligt i stoftet . 
Du behöver väl inte filma det ? 
Det var anledningen till att jag gick med på fyra . 
Du har helt fel synsätt på det . 
Du tjänar fyra miljoner pund på att medverka i filmen . 
Det är en miljon i minuten . 
Du blir världens bäst betalda skådis . 
Du borde fira , inte förhandla . 
Du , kompis ... - Det där kan förfölja mig för evigt . - Rör mig inte . 
Jag är inte din kompis . 
Det ska du ha klart för dig . 
Idag arbetar du för mig . 
Jag regisserar och du uppträder . 
Jag vill ha valuta för mina jävla pengar . 
Kom igen , Freddy . Det är bara en sång . Gör det bara . 
Dräkten . Uppträdandet . Kör . 
Jag ska bara gå och förbereda mig . 
Vill ni ha vargen i hönshuset ? 
Höna . Hö ... 
Du är en jävla Liverpool-tönt . 
Okej ! Nu kör vi . 
Var ska jag stå ? 
Ska du inte ta fram kameran ? 
Det funkar inte så . 
Du ska dansa . Sen avgör jag om uppträdandet är inspelningsvärdigt . 
Vet du varför du bär hönsdräkt ? 
För att förödmjuka mig inför hela jävla världen ? Det är inte en örndräkt av en anledning . Örnar dansar inte . De svävar fram . Genom luften . 
Men hönan är längst ner i näringskedjan . 
Du är en höna , eller hur ? 
Du kunde inte betala din skuld utan andras hjälp . 
Men du kan göra bot . 
Min bror gillar botgöring . 
Och en del av pengarna är hans . 
Han ser dansen som en liknelse . 
Just därför kan du inte bara låtsas vara en höna . Du måste vara en höna . 
Förstår du ? 
Botemedlet finns i giftet . 
- Kom igen . Visa oss din höna . 
- Okej . 
- Sätt igång . - Jaja ! 
Nej . Vad fan är det där ? 
Vad fan är det där för skithöna ? 
Kom igen ! Bli en jävla höna ! 
- Jävla sprätt . 
- Vagga som en höna ! 
Och lätet . 
Nej , det suger ! 
Rör på halsen . 
- Var en höna ! 
- Det är jag ju ! 
Du ska vara en höna . 
Du ska känna det . 
Du ska förvandlas till en höna . 
Det ska inte finnas nåt mänskligt kvar i dig . 
Jag vill bara se fågeln . 
Så kom igen . 
Få se . 
Vad gör du ? En höna går inte så . 
- Picka ! Lägg en äggjävel ! - Jag pickar ju ! 
- Jag pickar ! - Gå upp på soffan och flyg . 
- Jag är ett kukhuvud ! 
- Var en höna ! 
- Jag kan inte flyga ! 
- Var en jävla höna ! Kom hit ! 
Kom igen ! 
Titta , här finns korn . 
Picka på kornen ! Kom hit ! Och en mask . 
Ät upp masken , din jävla höna ! 
Kom hit ! Det är en mask här . En mask ! 
Picka på kornen ! Kom igen ! Picka på kornen ! Jag pickar ju , för fan ! 
Susie , vi måste stoppa det . 
Lägg dig inte i . 
Ät upp den jävla masken ! Ät upp den ! 
Ät upp masken , din jävla höna ! 
Tommy ! Det räcker nu ! 
Dra åt helvete ! 
Lägg dig inte i ! Annars ska jag ha mina åtta miljoner ! 
Kan du inte bara filma det så vi blir klara ? 
Han måste komma upp i hastighet först . 
Han måste bli en höna . 
Din jävel ! 
Kom igen ! Bli en höna ! 
Jag ... Jag måste gå på toa . 
Gå då , för fan ! 
Rappa på ! 
Hej , Tommy . Vem är det som är hönan nu ? 
- Freddy ! 
- Dra åt helvete ! 
Skjuten i pannan Som det kukhuvud han var Lian , lian , lej Lite pang-pang här Och lite pang-pang där En döing här , en döing där En döings hjärna överallt Nu har jag skjutit skallen av nån Lian , lian , lej ... 
