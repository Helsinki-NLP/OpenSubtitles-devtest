... förhållandena förvärras ... Varför svarar ni inte ? Det är flammor ... Eld ! Eld ! Kapseln har fattat eld . 
Tjugoett ... Tjugoett ... Trettio ... fyrtio ... fyrtiotvå ... Det är flammor ... 
Kan vi öka värmen lite ? 
Den är trasig , gumman . Svep in dig . 
Mamma ? Vad säger hon ? 
Hon säger att världen är uppochner . 
När kommer pappa ? 
Mamma ? 
Vad har hänt med pappa ? 
Stäng dörren , gumman . 
Åh , det är iskallt . 
Kom , jag ska tända brasan . 
Kan du berätta en saga ? 
- Jag kan läsa för dig . - Den på iPaden . 
Om rymden . Den är min favorit . 
Hej , jag heter Johanna . Jag är astronaut . Och jag arbetar för Europeiska rymdbyrån . Jag bor på den internationella rymdstationen . Jag ska vara här uppe i ett helt år , och jag har en väldigt speciell nattsaga . Den heter " Den lilla raketflickan " . 
- Vill du att jag läser den ? - Ja . 
Den lyder så här . " Uppe och ute i rymden är det väldigt kallt . 
Stjärnorna rör sig snabbt och solen brinner het bara för att hålla sig varm . 
Uppe och ute i rymden är det tyst . 
Men det värsta med rymden är att det kan vara väldigt , väldigt ensamt . " 
KÖLN - TYSKLAND Alice ? Vi åker om en kvart . 
Jag kommer . 
Avvakta . 
- Jag är klar att åka . - Okej . Hälsa . 
Kontrollcentret kopplar er nu . 
GEMENSAMT ÄGD AV NASA , ROSKOSMOS ( RYSSLAND ) , EUROPEISKA RYMDBYRÅN ( ESA ) , KANADA OCH JAPAN . God morgon , älskling . Har du borstat dina tänder ? Ja . Hur många minuter ? Tre minuter . 
Bra , för vi gör alltid tre minuter . 
Ska du på din rymdpromenad i dag ? 
Men du , du behöver inte vara orolig , baby . Det kommer gå så bra . 
Jag vet . 
Vill du säga god morgon till Yaz ? 
- Hej , Alice . God morgon . - Hej , Yaz . 
Är du nervös ? 
Bara lite . 
Vill du titta på salladen ? Den ser lite piggare ut , tycker jag . 
Den har liksom vaknat till lite . 
Vad tycker du ? 
- Är det inte magiskt ? 
- Wow , snyggt . 
Men jag låter nog - nån annan prova den först . - Ja . Jag är orolig att den förvandlar mig till en alien . 
Vi måste viska . Varför då ? 
För att de gör nåt väldigt pillrigt inne i CAL . 
Hej , Alice . 
Hej , Paul . 
Din mammas stora dag i dag . 
RPL . CAL-data : kärnsignalerna gröna , magneterna inriktade , 25,5 . 
- Uppfattat , fas sex . - Uppfattat . 
Kärntemperatur : minus 203 grader . RAKETDRIFTSLABORATORIET PASADENA , KALIFORNIEN Finjustera lasrarna . Kom igen . 
Vad gör den ? 
Den söker efter ett nytt materietillstånd . 
Vad betyder det ? 
Vet inte . 
Åttiofyra dagar tills du är hemma . Bara 84 . 
Jag längtar . 
Jag saknar dig så mycket . 
Jag saknar dig också , mamma . 
Tar du det försiktigt där ute ? Alltid . 
Få se om jag kan se dig . 
- Wow . - Titta . Där är du . Ser du ? 
- Vi är redo . - Då så . 
Lycka till , unge man . 
Lycka till , befälhavaren . 
Jag har haft turen med mig hittills . 
Hej , Alice . Vinka till dig själv . 
Sätt igång . 
Stationen , RPL , hör ni mig ? Få tillbaka dem . Vi är mitt uppe i nåt . 
Mamma ? Är du där ? 
Är allt okej ? 
Hon är borta . 
Rymdskrot ! Skrovet perforerat ! 
Mamma ? 
Houston , det här är Stationen . Hör ni mig ? 
Houston , det här är Stationen . Hör ni ? 
- Kontrollcentrum , lås dörrarna . - ... inte aktiverat . 
NASA : S KONTROLLCENTRUM Stationen , Houston på rymd-till-mark 1 , ni har en trycksänkning . 
Alla kanaler är öppna . 
Besättningen samlas i evakueringskapsel Sojuz 1 . 
Förbered evakuering . Verkställ krisrespons . 
Houston , brand och dimma i Zarja . 
- Stäng ner . - Ilja ! 
Jo , ta dig omedelbart till närmaste evakueringskapsel Sojuz 1 . 
Houston , det finns en brand mellan oss och Sojuz 1 . 
Samlas i Rassvet istället . 
Jo , jag kommer inte igenom ! 
Ilja , vi måste ta oss till evakueringskapseln ! 
Uppfattat . 
Vad fan träffades vi av ? Nåt träffade oss ! 
Ta dig igenom nu ! 
Jag är ute . 
Håll i mig ! 
Jag stänger luckan . 
Stationen , ni måste kväva branden . 
Uppfattat ! Fixar det ! 
Stänger av lufttryckssystemet i Zvezda . Nåt kolliderade med oss . 
- Är ni okej ? 
- Lucka säkrad . 
Besättning , upprop . 
Ericsson . 
Andrejev . 
- Brostin . 
- Suri . 
- Lancaster ? 
- Jag sitter fast . 
Luften är ren . 
Ericsson , Brostin , luften är ren . Hjälp befälhavare Lancaster . 
Uppfattat . 
Andrejev , Suri , kolla systemen och livsuppehållande . 
- Ska bli . 
- Kollar . 
Houston , vi förlorar syre . - Jag hör det . 
- Stationen , uppfattat . 
Paul ? Hur mår du ? 
- Jag sitter fast . 
- Han är fastkilad . 
- Han blockerar trycksänkningsreglaget . 
- Vi måste lägga förband här . - Sätt tryck mot pulsådern . - Jag fixar det . 
- Houston , Paul är skadad . 
- Uppfattat . 
Hans vänstra arm är krossad under ställ fyra . Han blöder kraftigt . 
Vad är statusen på systemen ? 
Ilja , vad är statusen ? 
Strömavbrott i 55 % av Zvezda och Quest . 
Tryckförlust i Harmony , Columbus . 
Jo du har ansvaret nu . 
Vi måste ge honom syrgas . - Uppfattat . 
- Sätt fart . 
Besättning , utvärdera evakueringskapselns livsduglighet . 
Ni signalerar allvarlig syre - och tryckförlust över hela ISS . 
Uppfattat . Ilja ? 
Paul , håll dig vaken . Audrey , du måste förbereda Paul för omedelbar evakuering . 
Andas . 
- Hör du mig ? - Han klarar inte en evakuering . 
Jo , elfel i kapseln Sojuz 1 . 
Signalerar 95 % elfel . 
Sojuz 2 funktionsduglig . Sojuz 1 skadad . 
Det finns bara tre platser i Sojuz 2 . Vi kan bara evakuera tre av oss . 
Svåra skador på alla livsuppehållande och övriga system . 
Avvakta . Ni kan i nuläget inte skjuta upp Sojuz 1 . 
Pumpa . 
Kan vi inte flytta honom , så måste vi amputera armen . Jag är ledsen , Paul . - Jo ... 
- Du kommer att klara dig . 
Jo ? Ilja ? Ni hade en rymdpromenad på schemat denna morgon . 
Ni måste fullfölja den för att laga det livsuppehållande systemet och skadorna på Sojuz 1 . 
Jag vill vakna igen . Okej . Han är medvetslös . Vad gör vi med Paul ? 
Jo , Audrey kan ta hand om Paul . Uppfattat . 
Ni måste undersöka skadorna på evakueringskapseln i Sojuz 1 . Laga livsuppehållande system och elfel . - Uppfattat . 
- Sen kan vi få hem er . 
Framme . 
Okej , kom . Usch . Vi får inte båda bli sena . 
Om ni är uppmärksamma , så var vi sex sekunder in i lasersändningen när olyckan inträffade . 
CAL skulle ha tagit emot information inom två miljondelars sekund . 
Håll tempen under minus 120 grader och ordna en räddningsplan . 
Befälhavaren , vi får en signal från CAL . En sändning går fram . 
Irena Lysenko , Roskosmos . 
Befälhavare Henry Caldera , - vetenskaplig chefskonsult ... - Henry . ... på Raketdriftslaboratoriet . 
- Titta . - Michaela Moyone , NASA:s kontrollcentrum . 
- Herregud . - Frederic Duverger , chef för Europeiska rymdbyrån . 
- Vi hade en kraftig kollision ... - Kom . Har du sett det här ? - ... på ISS ... - Herrejävlar . ... och vi måste diskutera full evakuering . 
Alice , hej , kom här . 
Okej , sätt er på era platser , allihop . 
- God morgon . - God morgon . 
Är du okej , Wendy ? 
Jag hade mardrömmar . 
Jo , Ilja , ert mål är att bedöma skadorna på de elektriska och livsuppehållande systemen . Förstått . 
Okej , Jo . Du har klartecken för lucköppning . 
Uppfattat . 
Luckan är öppen och säkrad . - Jag är på väg ut . 
- Jag är precis bakom dig , Jo . 
Jo , Ilja , jag lämnar över er till Roskosmos kontrollcentrum under er rymdpromenad . 
Lycka till . 
Uppfattat . Förstått . 
Vi instruerar . Låt oss få det åtgärdat . 
ROSKOSMOS KONTROLLCENTRUM BAJKONUR , KAZAKSTAN Okej , vi är båda igenom luckan . Det kommer att vara mörkt i ytterligare cirka 20 minuter . 
Uppfattat . 
Jo , Sojuz 1-kapseln signalerar fullständigt strömavbrott . 
Ni måste laga elkablarna på Unity . 
Uppfattat . 
Ilja , bege dig ner för att undersöka evakueringskapsel Sojuz 2 . 
Uppfattat . 
Ovanför Nauka , cirka åtta meter . 
En del ytliga skador . 
Men Sojuz 2 ser ut att vara mer eller mindre intakt . 
Houston , Stationen här . Operation genomförd på Paul . 
Uppfattat . 
Stationens livsuppehållande system är nere på 30 % . 
ESA , ni kan inte nog betona vikten av detta experiment . 
Vi fick en signal . En dubbelkvantumsignal . Det är oerhört betydelsefullt . KÖLN , TYSKLAND Vi förstår betydelsen , RPL , men vi kan inte prioritera NASA-experiment över en evakuering . 
Läxa inte upp mig om evakueringen , Frederic . 
Jag har hållit på med det här i 50 år . 
Om vi överger ISS i det rådande politiska klimatet , kommer vi aldrig att återvända . 
NASA , vetenskapen är inte viktigare än människorna . 
Vi driver inget djävla dagis där uppe . 
Vi har hittat ett nytt materietillstånd som bara kan existera i tyngdlöshet . 
Vad felet än är där uppe , så kan det åtgärdas . 
Vi har allvarliga kollisionsskador på strömförsörjningen . 
Syresystemet , yttre elkablar avskurna från den här sidan . 
Kan ej kopplas in igen . 
Skador irreparabla . 
Houston , direktiv , tack . 
Paul håller på att få hjärtstopp . 
Inleder HLR . 
Ett och två och tre och fyr och fem och sex ... Avbryt rymdpromenad . Avbryt rymdpromenad . 
Förbered Sojuz 2 för omedelbart återinträde . 
EVA och Houston , bortse från den ordern . - Vi är inte överens . - RPL . Houston , håll den här kretsen öppen . 
Jag tillåter inte att vi fattar det beslutet förrän vi har kalkylerna för att rädda CAL-experimentet . 
Oenig . Nu avslutar vi samtalet och får ner dem därifrån . 
Sergej . Fortsätt med rymdpromenaden . 
Jo , sjukvårdsteamet tar hand om Paul . Fortsätt med rymdpromenaden . 
Uppfattat . 
Håll mig uppdaterad . 
Vart ska jag nu ? 
Skicka henne till truss . De måste åtgärda sekundära livsuppehållande system . 
Vad är problemet ? Jo , vi kan inte se vad du ser . 
Den lyser rött . 
Det är nåt fel . Tyvärr . Vi har inga kameror igång bortanför Unity . 
Hon måste fortsätta . 
Okej . En minut till soluppgången . 
27 , 28 , 29 , 30 . 
Solljus om fem , fyra , tre , två , ett . Jo , du måste till truss för att laga sekundära livsuppehållande system , annars har besättningen varken ström eller syre för att reparera Sojuz 1 . Uppfattat . 
Vi har inga kameror på truss . Alla är avstängda . 
Vi flyger i blindo från och med nu . Okej . På väg till de sekundära livsuppehållande systemen . 
28 , 29 , 30 . 
- Sluta . - Undan . 
- Börja . 
Truss kommer inom synfält . 
Hämta amiodaron . 
21 , 22 , 23 , 24 , 25 , 26 , 27 . 
Vad som än träffade oss totalförstörde de sekundära livsuppehållande systemen . 
Det här var en kraftig kollision . 
Ett och två och tre och fyr ... - Kan du se vad som orsakade den ? 
Jag närmar mig . 
Ser ut att vara en ... reva på kanske 50 centimeter . 
Nåt är intrasslat i ... i truss . 
Ilja , uppfattar du ? 
Jag är nästan där . 
Jo , bekräfta vad du ser , tack . 
Det är orange tyg . 
Jag tror jag måste titta ovanifrån . 
Kom tillbaka . Helvete . Det är en kropp . 
Jo , vänligen bekräfta . 
Jo , svara . 
Ilja , vi behöver kameror på Ericsson . 
Jo ! Jag kommer ! 
Kolla min syrgas . 
Kom igen , Jo . 
Jag har dig . 
Hon är i säkerhet . 
Fråga om han ser nåt . 
Andrejev , ser du nåt ? 
Nej . 
Det var en kvinna . CCCP . Sovjet . 
Jag såg en död kvinnlig kosmonaut . 
Kom igen ! Kom igen , jag ger inte upp ! 
Houston , TsUP Paul är död . 
Jag upprepar , befälhavare Lancaster är död . 
Jag ... Jag är ledsen att behöva vidarebefordra det här . Stationen rapporterar att befälhavare Lancaster har avlidit . 
Han har avlidit till följd av hjärtstopp . 
Farväl , Paul . 
Sojuz 2 , förberedelser för avdockning slutförda . 
Utträdesparametrar upplänkade . Anhöriga på väg till Bajkonur . 
Det gör fan ingen nytta om vi alla är döda . 
Ta det lugnt . 
Vi har ett reparationsschema för Sojuz 1 . 
Tre av er åker nu i Sojuz 2 . Den kvarvarande besättningsmedlemmen lagar elskador i Sojuz 1 med hjälp av 606-batterier från den ryska befälsmodulen . 
Sen har Sojuz 1 klartecken att återvända . 
Varför åker inte två nu i Sojuz 2 och två stannar och reparerar Sojuz 1 ? 
Det livsuppehållande systemet kan bara hålla en person vid liv . 
Så , Ilja , Yaz Audrey , ni kom upp i Sojuz 2 . 
Jo , jag stannar . 
Nej , du är befälhavare på Sojuz . 
Du ser till att få hem dem . 
Det är en order . 
Och Alice ? 
Vi har alla familjer . 
Lite klibbigt , eller hur ? 
Vet du , Luka , vi kan väl bara ta av vingarna och ... Eller vi kanske bara ska börja om ? 
Kommer hon tillbaka ? 
Jag hoppas det . 
Varför säger du inte ja ? 
Jag vill inte ljuga . 
Lyssna , stumpan . 
Mamma har alla möjligheter att komma tillbaka , men det är knepigt . 
Ingen har nånsin inte kommit tillbaka från rymden . Inte från en ESA-flygning . 
Jag måste berätta en sak . 
Det är upprörande . 
Tyvärr har Wendys pappa dött . 
Vad ska vi göra med våra cyklar ? 
Vi lämnade våra cyklar . 
Varaktighet av SKD-bränning , två minuter och 57 sekunder . 
- Inträdesvinkel , 95 grader . - Redo för avfärd ? 
- Parametrarna är inställda . 
- Redo för avfärd . 
Nåt du vill att vi ska säga ? 
Till dem där hemma ? 
Om jag inte kommer tillbaka , är du snäll och tar hand om Magnus och Alice ? 
Lutar station . 
Raketmotorer testade . 
Full styrka . Lossa . 
Uppfattat . 
Bultar apterade . 
Tänd raketmotor , KDU-motorer om tre , två , ett . Mekanisk frånkoppling . 
Jag ser separation . 
Går in i inflygningsbana . 
Tid till landning : tre timmar och 27 minuter . 
Om Gud så vill . 
Jo , du ska fylla Sojuz 1 med proviant för 24 timmar . 
Hur mycket livsuppehållande har jag ? 
Hur mycket syre ? 
Cirka 19 timmar . 
- Lyssna . - Sätt dig längst bak . 
- Jag ber om ursäkt än en gång . - Ja . Herregud . Jag är hemskt ledsen . Wendy , du kan väl sätta dig hos Alice ? 
Jag är så ledsen , Frida . 
Vill du ha min kanin ? 
Sojuz 1 är skadad . 
Den har andningsbar atmosfär men inte nog med ström för att ta dig hem . 
När du har fyllt Sojuz 1 med proviant , måste du avlägsna de döda batterierna och ersätta dem med 606-batterierna uppe i Zvezda . 
Du kommer att ha syre och ström i ISS var 45:e minut för reparationer . 
Uppfattat . 
Jo , din familj är på väg . 
Du kan prata med dem när det blir ljust igen . Toppen . 
Stäng huvudluckan . 
- Trycksätt . 
- Uppfattat . 
Vänta . 
- Jag kommer strax . - Jo , ISS har bara solkraft nog för belysning och livsuppehållande . 
Du har en och en halv minut . 
Kvällningen kommer . Du kommer inte att kunna trycksätta . 
Jag måste bara hämta en sak . Jag hinner i tid . 
Jo , under natten kommer du bara att ha syre i Sojuz 1 . 
Jag vet . 
- Jo . 
- Hälsa Alice att jag tar hennes halsband . 
- Jo , 20 sekunder . 
Mamma älskar henne . Det betyder att jag klarar mig . 
Jag kommer hem till henne och pappa . 
Lova att hälsa dem det . Tio , nio ... - Lova att säga det . - ... åtta sju , sex ... Sergej , lovar du ? 
Om du inte lovar , kommer jag bara att sitta här och tjura . 
- Vi ska framföra det . 
- Tack . 
Så , det här är proceduren varje omlopp : Fyrtiofem minuter i dagsljus , 45 minuter i mörker . 
Pausar kommunikation . Åter i dagsljus om fyrtio ... 
För protokollet , och jag vet hur historiskt osannolikt det är , det här är min skildring av vad som träffade solpanelerna . 
Liket av en kvinna i sovjetisk rymddräkt . 
Ska vi leta upp mamma , Alice ? 
Åh , min älskling . 
God morgon , Stationen . God morgon , Jo . God morgon , Sergej . 
- Du är alltid så munter . 
- Tack , Jo . 
Vi har cirka 17 timmar och 49 minuter . 
Låt oss leta upp batterierna . 
Det gör vi . Jag vill komma hem . 
Batterierna byggdes inte för att flyttas , men bör vara åtkomliga . Förstått . 
Det kommer att ta längre tid än vi trodde . 
SKD om minus 20 . 
Tänder raketmotor om fem , fyra , tre , två , en . Separation fullbordad . 
Irena , du är ansvarig för den här jäkla evakueringen . 
Jag skickade dig en plan . 
Jag vill att Ericsson tar med sig CAL tillbaka . 
Henry , jag instruerade dem att lämna din maskin . 
Varför i hela friden då ? 
Såvitt jag vet , orsakade den olyckan . 
Irena , det finns nåt inneslutet i de sex sekunder den var i drift som kan förändra allt . 
För dig , för mig , min bror . 
Den fungerade . Vi måste få tillbaka den . 
Vi får inte fler chanser . 
Skicka räddningsplanen , snälla . 
Sojuz 2 , bekräfta parametrar för omloppsutträde . 
Bekräftat . Träder in i atmosfären . 
Kapseln har återinträtt i atmosfären . 
Skicka räddningsplanen för CAL . 
Ja ? Jag går just av planet . 
Jag går direkt till kontrollcentret . Vad är hennes status ? 
Okej . Ja . Hej då . 
Det blir snart natt hos henne . Om vi skyndar oss , kan ni prata med henne . 
- Bra . - Ja ? 
Spänn åt alla era remmar hårt när ni är under G. 
Försök hålla era luftvägar öppna genom att luta huvudet bakåt . 
Radioavbrott . 
TsUP , har ni uppfattat ? 
Vi hör dig , Ilja . Klart och tydligt . 
Skönt att höra era röster . 
Sojuz 2 utlöser fallskärm , går in i kontrollerad landning . 
Jo . Goda nyheter . Sojuz 2 har landat . 
Uppfattat . Toppen . 
Jo , vi skickar några ritningar . 
RPL har begärt att du räddar ett av deras experiment . 
- Vilket experiment ? 
- CAL:s datakärna i Destiny . 
Det känner jag inte till . Vet inte om jag hinner . 
Det är ett NASA-experiment . Äventyra inte din säkerhet . 
Är min familj där ? 
De är på väg . 
- Tio minuter till kvällning . - Uppfattat . 
Jag vet att du och mamma hade problem . 
Men jag vill att ni ska vara vänner vad som än händer . 
Din familj är här och kommer för att prata med dig . 
Jag vill gärna prata med dem också . 
Underbart . Vi ordnar det . 
Uppfattat . 
Låt oss fixa batteriet innan kvällningen . Det gör vi . 
Din familj kommer in nu . Uppfattat ... Stationen , det här är TsUP . 
TsUP , Stationen här , kom . 
TsUP , Stationen här , kom . 
Vad händer ? Pappa , vad händer ? 
Hallå , Stationen här . Är min familj där ? 
Jag ska fråga vad som hänt . Stanna här en sekund . 
Ursäkta ? Hallå ? Ursäkta ? 
Vad händer ? 
Snälla , svara . 
Alice . Kom tillbaka . Alice ! 
Va ... 
Var har du varit ? 
