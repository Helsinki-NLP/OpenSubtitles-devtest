Frukost , ungar ! 
Lugn . Ingen brådska . 
Det finns gott om pannkakor . 
- Tack , mamma . Älskar dig . 
- Tack , mamma . Älskar dig . 
Jag älskar er också . 
Och jag , då ? 
- Dig med , pappa . - Dig med , pappa . 
Raring , har du varit till frissan ? 
Du är jättefin . 
Bara en liten putsning . 
Vi har slut på Honey Pops . 
Ursäkta ? 
Vi har slut på Honey Pops . 
Carlotta ? 
Honey Pops . 
Vi har slut på Honey Pops . 
Carlotta ? 
Carlotta ! 
Honey Pops ? 
Och vad ska jag göra åt den saken ? 
Mår du bra ? 
Du ser trött ut . 
Jadå . Jag mår bra . 
Jag ser alla dessa människor som lever sina liv som om inget hänt ... Dedo , vi har hållit på i flera veckor nu . 
Vi är inte närmare att hitta Wanda , känns det som . 
Intendent Rauch avspisar mig . Så polisen är tydligen inte närmare lösningen än vi . 
Det är bara en tidsfråga . 
Vi får ett genombrott snart , det känner jag på mig . 
Ole föreslog att pröva med en drönare med värmekamera . 
Ska vi köpa en ? Vad tycker du ? 
Värt att chansa ? 
Ta ledigt idag , vetja . Få lite frisk luft , ta en simtur . 
Så fortsätter vi imorgon . 
Jag fortsätter bevaka ett tag till . 
Då känner jag att jag gör nånting . 
Som du vill . 
Jag går och gör en smörgås . 
För cirka hundra år sen definierade schweizaren C.G. Jung synkronicitet som händelser som verkar inträffa samtidigt av en slump men som ändå hänger samman och bara kan förstås tillsammans . 
Ärligt talat var han lite överdriven . 20 M - ANDRA AVFARTEN 
Jag menar , har ni nånsin tänkt på hur många saker som måste hända tillsammans , samtidigt , för att till slut allt ska bli precis som det blir ? 
Tänk om bara en enda detalj var annorlunda ? 
Ert liv skulle ta en helt annan bana . 
Som när min mamma tyckte att det var en bra idé att vår granne Karin skulle frisera mig , och så gav hon mig en jätteful lugg som gjorde hela skolåret i trean till ett helvete . 
Ödet kan vara ett riktigt rövhål ibland . DAG 96 Wanda åker hemifrån . 
Hennes mobil återfinns på kaféet . 
Här kastas hennes T-shirt i containern , och här syns hon i Lenkas Instagraminlägg . 
Mobildata från Lenkas mobil visar att hon stannade här , här , här , här och här , innan hon tydligen körde utan uppehåll hela vägen tillbaka till Tjeckien tills hon körde nedför ett stup . 
Hon kanske somnade vid ratten ? Trött av långkörningen . 
Det liknar nästan en mus . 
Nosen , öronen och svansen . 
Så fotot vid statyn är Lenkas sista inlägg . 
Och den dessförinnan var här . 
LENKA-UNDERSÖKER # INVESTIGATIVEINFLUENCER Hejsan . 
Hittade ni den skyldiga ? 
Den som åt upp era fåglar . 
Just det , fåglarna . 
Ja . 
Vi tror att det är en grävling . 
En grävling ! 
Vilket majestätiskt djur . 
Men de brukar inte ta fåglar . 
Inte ? 
Men den här jäkeln gör det . 
Just det . 
Hursomhelst tänkte vi genomsöka skogen för att hitta grytet . 
Min son talade om drönare med värmekamera . 
Jag har precis vad ni söker . 
En grävling ? 
Allvarligt ? 
Lucie , smyger du dig på mig ? 
Du vet att jag inte tycker om det . 
- Är allt okej ? - Jadå . 
Ja ? 
Förlåt , vännen . Ursäkta mig ett ögonblick . 
Vad är det ? 
Det passar inte så bra ... Hej , det är jag . 
Jag försökte prata med mamma igen , men hon är för upptagen . 
Jag börjar bli lite rädd , men det är förmodligen ingen fara . 
Jag menar , Lina hade inte mens på två veckor , men det var för att Merkurius var på bakåtgående . 
Ring tillbaka , snälla . 
Oj , alltså . 
- Varsågod . 
- Tack . 
Har du nånsin krossat en mans hjärta ? 
Harald ! Vad har vi sagt om att skrämma bort kunder ? 
Förlåt . 
Hans fru har kommit på ett boende för dementa . 
Åh , jag beklagar . 
Och hans flickvän lämnade honom . 
- Allt väl , Harald ? - Jadå . 
Vad önskas ? 
Jag utreder försvinnandet av en ung kvinna . 
Wanda Klatt . 
Ja . Jag känner familjen . 
Det är hemskt . 
Anita ! 
Harald ! 
Jag menar en annan kvinna . Jaha . 
Henne känner jag inte . 
- Vem är hon ? 
- En influencer från Tjeckien . 
Såna tillhör inte vårt vanliga klientel . 
Hon var här Nuppelwocken-kvällen . 
Det kommer massor av människor hit då . 
Det är nog vår bästa kväll på hela året , med paraden och fotbollen ... 
- Varför söker du henne ? 
- Hon är död . - Död ? 
- Hon dog i en bilolycka . 
Antas det . 
- Vid tjeckiska gränsen . - Ja . 
- Knappt ett dygn efter att hon var här . - Herregud . 
Jaha , ja . 
Nej . 
Nej . Henne minns jag inte . Beklagar . 
Okej . 
- Ifall du kommer på nåt . - Så ringer jag . 
- Hej då . - Hej då . 
- Harald , igen ? Allvarligt ? 
- Anita . Ja , Anita . 
- Här . 
- Vad tar du dig till ? 
Vadå ? 
Idag är leveransdag . 
Sista avbetalningen görs idag . 
Inte här . 
Följ med mig . 
Hej . Vad önskas ? 
En ananasjuice med tequila , tack . 
Men ananasjuicen måste vara färsk . 
Okej , jag tar en sån där . 
Tjusig utstyrsel . 
Vad föreställer du ? En fågelskrämma ? 
Jag föreställer Nuppelwocken . 
Ikväll är Nuppelwocken-kvällen . 
Wuppelnocken ? 
Nuppelwocken ! 
Puppen-Dockel ? 
- Nuppelwocken . 
- Jag förstår inte vad du säger . 
Det är en gammal legend . 
Se där . 
Det är Nuppelwocken , ett monster som lever i skogen och vart hundrade år kommer hit och rövar bort den skönaste jungfrun . 
Coolt . 
Så jag får passa mig . 
Gör det du . 
- Önskas nåt mer ? - Ja , visst . 
Vet du vad en myrkott är ? 
- Va ? 
- De är så söta . 
Men fler än en miljon myrkottar infångades olagligt bara förra året . 
Sluta filma , tack . 
Jag försöker spåra upp hjärnan bakom Europas största liga som smugglar vilda djur . 
Jag bad dig snällt att sluta filma . 
Han kallar sig King . 
- Hon sa ju åt dig . - Hallå . 
Om du rör mina grejer igen , Voldemort , får du pepparsprej i snoken . 
Hör på ... Jag har aldrig hört talas om nån " King " . Så drick upp och ge dig iväg . 
- Har du inte ? 
- Nix . 
Märkligt . 
För han gör sina affärer här . 
Black Souk . 
Vet du vad det är ? 
En marknadsplats på mörka webben . 
Ett misstag många människor gör är att tro att mörka webben är totalt anonym . 
Men det gör dem sårbara . 
Vänta här . 
Vad är det ? 
Glo inte på mig så där . 
Jag har 125 000 följare . 
Jag kan skicka min trollarmé på dig . 
King vill prata med dig . 
Skriv din kontaktinfo . 
X , TikTok eller Insta ? 
Ditt telefonnummer . 
Okej , gamling . 
Förresten smakar ölen skit . 
Ja , det är jag . Du måste komma genast . 
Nej , tack . 
Det är enda bussen som går härifrån . 
Jag tar nästa . Tack . 
Nästa kommer om en timme . 
Jag väntar , tack . 
- Vill du prova ? 
- Det är nog ingen bra idé . 
Få se vad den kan göra . 
Och hur är det med dig ? 
Mår du bra ? 
Det har varit lite galet på sistone . 
Att mista Wanda så där plötsligt . Utan förklaring . Det påverkar en . 
Det får en att inse hur små vi är i detta jättestora , kaotiska universum . 
Som små möss som springer omkring på järnvägsspåret . 
Omedvetna om att de kan krossas när som helst . 
Men när man får se världen så där , kan man inte glömma det . 
Hur slutar det ? 
Vad menar du ? 
Tänk om vi inte hittar henne ? 
Vi ska hitta henne . 
Vi måste . 
Okej , få se nu . 
Var är vi ? 
Det där ser bekant ut . 
Det är det nya kebabstället som just öppnat . 
Ska vi äta lunch där efteråt ? 
En klasskamrat gick dit . 
Var kebaben bra ? 
Han sket på sig på bion senare . 
Hamburgare , alltså ? 
Så , härifrån går man norrut till gatukorsningen . 
Man följer huvudleden till rondellen . 
Förbi hyreshusen . 
Fortsätt , fortsätt . 
Och så stanna vid hörnet . Stopp . 
Precis där . 
Det är vår startpunkt . 
Där allt började . 
Containern där de fann Wandas T-shirt . 
Ta upp den så högt det går nu . 
INSAMLINGSCONTAINER Vi har kollat alla de här . 
De där också . De enda som återstår är de här och husen vid skogskanten . 
Åh , Wanda , vännen , vi vet att du finns där nånstans . 
Ge oss ett tecken . 
Wanda ! 
- Wanda ! 
- Wanda ! 
- Var är du ? 
- Wanda ! 
- Hej , Lucie . 
- Hej . 
Vi går i skolan ihop . 
Alla är ungefär likadana . 
Jag skulle ta den här . 
Den finns i tvåpack . Och den är superenkel . 
Jag köper för en vän . 
Hälsa din vän att hon inte behöver vara generad . 
Nästan varenda kvinna har gått igenom samma sak nån gång . 
Men vi pratar inte om det . 
Jag pratade aldrig om det med min dotter heller . 
Jag trodde väl att om jag inte pratade om det , så skulle det inte hända . 
Rätt dumt , eller hur ? 
När jag försöker prata med mamma om det har hon inte tid . 
Lucie , tro mig , hon har alltid tid för att prata om det här . 
Hur vet du vad jag heter ? 
Du går i samma skola som mina barn . 
Jag ... Jag är Oles och Wandas mamma . 
Du verkade bekant . Ja . 
Jag är ledsen för det här med Wanda . 
Hon var cool . Hoppas hon kommer hem . 
Jag menade inte att ... Behöver du sätta dig ? 
Vi kan ta en kaffe eller nåt . 
Visst . Vi dricker kaffe . 
Oj , gott , va ? 
Gissa vem vi kan rekommendera Spicy Snacks till ? 
Morbror Rüdiger . 
Han skulle nog gilla det . 
Det var kul att hänga . 
Vi borde göra det oftare . 
Det är inte så lätt . 
Du och mamma är jämt upptagna med det här med Wanda . 
Men vi har alltid tid för dig också . 
Det vet du väl ? 
Ska du och mamma skiljas ? 
Va ? 
Nej . 
Varför tror du det ? 
Har mamma sagt nåt ? Nej , nej . 
Men hon är arg jämt , och du gör saker som retar upp henne . 
Kompis , jag försöker verkligen . 
Jag vet . 
Va ? Vad är det här ? 
Jäklar . 
Han hittade kameran . 
Inte bra . 
Polisen ? 
Nån har brutit sig in hos mig . 
Inte bra alls . 
- Ska vi ringa mamma ? - Nej . 
Vi grejar detta . Kom igen . 
Vi måste bara få bort kamerorna därifrån . 
Det var snällt av dig . 
Jag mår redan bättre . 
Jag vet inte riktigt vad det var . 
Det är okej . 
Jag fattar . 
Det måste vara tufft . 
Wanda går i klassen över mig , men jag minns henne . 
Hon var jämt så tjusig och rolig . 
Sån är hon . 
Jag mötte nån morgonen hon försvann . 
I skogen . 
Du är sen . 
Jag tog en omväg för att inte bli sedd . Hela stan är i farten idag . 
Men ingen såg dig väl ? 
Slappna av . 
Du är så paranoid . 
Jag kan mista jobbet . 
Du är 15 . 
Jag kan få fängelse . 
Ingen såg mig . 
Jag lovar . 
Och jag såg Wanda . 
Berättade du för polisen ? 
Varför inte ? 
Det här är viktigt . 
Förlåt . Jag är så ledsen . 
Jag vet att jag borde ha sagt nåt . 
Jag ville säga nåt , men jag ... Jag måste lova honom att inget säga . Vem fick dig att lova det ? 
Han är lärare . 
Okej . Jag förstår . 
Och jag antar att det är skälet till det här ? 
Åh , Lucie . 
- Lucie , Lucie ... 
- Säg inget till mamma , snälla . 
Okej . 
Jag ska inget säga till henne . 
Herr Hessel , det är polisen . 
Vad vill ni mig ? 
Hjälp ! 
Varför gör han sånt motstånd ? 
Inte bra . Inte bra alls . 
- Ta kamerorna . 
- Släpp , skitstövel ! 
Ni är ena riktiga fegisar . 
Ni ger er på fel kille . Jag har varit i armén . 
Varför slog du till honom så hårt ? 
Det var självförsvar . 
- Är han död ? 
Han ser inte ut att andas . 
Åh nej . 
Varför måste han skrika åt mig så där ? 
- Herregud . 
Vad har vi gjort ? 
- Vad gör vi nu ? 
... jag följer utredningen om Wanda på sociala medier . 
Massor av människor gör inlägg . 
Verkligen ? 
Har du hört talas om Mörka huset ? 
Mörka huset ? 
Ett hus på Forststraße . 
Det sista på vänster hand . 
Ingen går nånsin in och ingen kommer ut därifrån . 
Det har en hemsk grå färg , som ruttnande kött . 
Där finns skyltar med texten " Tillträde förbjudet " och " Argsint hund " . 
Men ingen har hört hundskall . 
En del säger att de som bor där hålls i skogen nattetid . 
De går bara ut i mörkret , vid fullmåne . 
Sökande efter nästa offer att uppsluka . 
- Vänta . 
- Det är bara en av teorierna . 
Andra tror att Wanda rymde för att bli med i Cirque du Soleil . 
Du vet , om du vill kan du kila in och ta provet nu . 
Jag är säker på att det är negativt . 
Men om inte , kan vi tillsammans räkna ut vad du ska göra . 
DAG 0 
King . Oj , du är inte vad jag väntade mig . 
Jag vet att du är en upptagen smugglare , så jag ska komma till saken . 
Antingen säger jag vad jag vet till polisen , eller så ger du mig en exklusiv anonym intervju . 
Jag har redan gjort en video som ligger låst och klar i mina utkast , klar att läggas ut . 
Frågan är , vill du att jag styr narrativet ? 
Va ? 
Allvarligt ? 
Okej , skicka plats , så kommer jag . 
Kom hit . 
Lucie , hör på . 
Du och den här mannen är nog ingen bra idé . 
Det finns väldigt bra killar i din egen ålder . 
Som min son , Ole . 
Jag är nog inte Oles typ . 
Försök inte med mig , kompis . 
Oj , alltså . 
Vi har alltså en död influencer och en försvunnen flicka . 
Kunde inte nån annan ha tagit hand om det här ? 
Vi har viktigare saker att göra . 
Herr Hessel . 
Ni ringde ? 
Det är Rauch från polisen . 
Öppna dörren , tack . 
- Tyst . 
Vad ska vi göra ? - Herr Hessel ? Är ni där ? 
Jag vet inte ... 
Vi tar bakdörren . 
Bra idé . 
Herr Hessel ? 
Var är skåpbilen ? 
Den stod ju här . 
Okej , herr Hessel . Vi kommer in . 
Vad ska vi göra ? 
Vi måste iväg . 
Sakta , mycket sakta . 
Spring ! 
Fan också . 
Tack för ... Du vet . 
Ingen orsak . 
Bara en sak . 
Morgonen du såg Wanda , åt vilket håll åkte hon ? 
Hon åkte åt det hållet . 
Men hon var ensam . 
Bra att veta . 
Tack . 
Lucie ? 
- Vad gör du här ? 
- Hej . 
Vi har träffats . 
Jag är Carlotta Klatt . 
Oles mamma ? 
- Och Wandas . 
- Herregud , javisst . 
Jag har sett dig vid skolevenemang . 
Du är potatissalladens drottning . 
Ja , Lucie ... Hon såg mig och ville uttrycka sin sympati . 
Jag visste inte att min dotter var så empatisk . 
Det har hon dolt från mig . 
Jag ville ha lite glass , bara . 
Vi kanske kan se en film tillsammans senare ? 
Jättegärna . 
Du kan väl gå in och välja en ? Jag kommer strax . 
Vi kan väl åka hem efteråt ? 
Jag ville bara säga att jag inte kan föreställa mig vad du går igenom . 
Om du vill ta en kopp kaffe eller bara nån att prata med , så bor jag strax intill . 
- Hemskt gärna . 
Tack så mycket . - Okej ? Bra . 
Skriv in ditt nummer , så sms:ar jag . 
Jösses . 
- En del kör som idioter . - Ja . 
Följer de efter oss ? 
Jag tror inte det . 
Ska jag svara ? 
Din mamma får aldrig veta det här , förstått ? 
Vilket då ? 
Att vi bröt oss in hos Hessel och slog till honom i ansiktet ? 
Eller att vi stal en skåpbil och flydde från snuten ? 
Herregud . 
Jag är inte dum . Klart att jag inget säger . 
Hon skulle slå ihjäl mig . 
- Det skulle hon . 
- Det skulle hon absolut . 
Sen få dig återupplivad på sjukhuset - så att hon kan döda dig igen . 
- Ja . 
Dig sätter hon i en internatskola i Schweiz där alla talar latin och klär sig som Harry Potter . 
Ta vänster här , tack . 
Stanna här . 
Okej , Utmärkt . 
Vi dumpar skåpbilen i skogen . 
Vad är det där ? 
FÖLJESEDEL LEVERERAS TILL : RÜDIGER SCHÄFER Rüdiger ? 
Va ? 
Pappa ! 
3 MISSADE SAMTAL CARLOTTA En hemlig övervakningskamera ? 
Just det . 
Dold i lampan i hallen . 
- Och det var två män . - Hej då . En kort och rund , och en mager . 
Med snabbmatpåsar över huvudet ? Just det . 
De bröt sig in och angrep mig . Slog mig medvetslös . 
När jag vaknade var både kameran och männen borta . 
Försvunna som genom ett trollslag , va ? 
Nu förstår jag allting . 
Det var så de visste om Margaret . 
Det var deras fel att Anita lämnade mig . 
Herr Hessel , minns ni att vi nästan stötte på varann häromdagen ? 
På Kapitän ? 
Var ni där länge till ? 
Fortsatte ni dricka ? 
Bara en tår på tand för att lindra sorgen . 
Anita är borta . 
Hon är borta . 
- Hon är borta . - Rauch här . 
Borta . 
Anita är borta . 
Fröken Rauch , det här är Carlotta Klatt . 
Jag vill bara berätta att nån såg Wanda . Dagen hon försvann , på väg in i skogen . 
Vad ? Hur vet ni det ? 
Jag talade med ett vittne . 
Vad för vittne ? 
- Det kan jag tyvärr inte berätta . - Ursäkta ? 
Det spelar ingen roll . 
Det här är ny information som ni inte hade . 
Fru Klatt , om informationen är trovärdig måste vittnet träda fram och uttala sig . 
Har ni redan undersökt Mörka huset ? 
- Vadå ? - Det stora , kusliga huset nära Forstplatz ? 
Det finns många , många teorier om det online . 
Några av dem är visserligen lite långsökta ... Jag stoppar er där , för jag har riktigt polisarbete att utföra . 
Men jag avråder från att söka efter Wanda på nätet . 
Ni hittar inget gott där . 
Adjö . 
- Dumma kossa . 
- Dumma kossa . 
Ole ! Snälla ! 
Ole ! 
Vakna ! 
Är du oskadd ? 
Ole . Hallå . Ole ! 
Är du oskadd ? 
Är du oskadd ? 
- Jadå . 
- Tack och lov . 
Förlåt mig . Jag vet inte vad som hände . 
- Mår du bra ? 
- Ingen fara , pappa . 
- Jag mår bra . 
- Herregud . 
Vi måste bort härifrån . Okej ? 
Oj , jäklar . 
Oj , jäklar . 
Herregud . 
Herregud . 
Pappa ? 
Varför finns det en bur inuti ? 
Ingen aning , och jag vill inte veta . 
Ge mig den där . 
Kom så sticker vi . 
Ole , kom nu ! 
- Mår du bra ? 
- Jadå . 
Har du ont nånstans ? 
Nej . 
Fan också . 
Har du kört vilse ? 
- Du är journalisten , va ? 
- Undersökande influencer . 
Samma som en journalist men med fler likes . 
Så du vill prata med King ? Ja . 
Följ med mig . 
Kom nu . 
Jag bits inte . 
Nej ! 
