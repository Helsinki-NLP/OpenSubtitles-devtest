Jag vet inte vad du hoppas kunna uppnå , Anna . 
Jag har försökt , den går inte att laga . 
Jaså ? 
Titta , du har fått tillbaka din vagn . 
Jösses . Jag hade fel igen . 
Vad skulle vår familj göra utan dig ? 
Din begåvning kommer att förändra världen . 
Men det är upp till dig hur du nyttjar den . 
Pappa ? 
Församlingen . 
- De ska väl inte ... 
- Gruvorna . De beslagtar dem . 
Gå ! Fort ! 
Magiker ! 
Perfekt . 
Pappa ? 
Anna ... Spring ! 
- Hur många själar ? - Över 500 döda . Åttahundra skadade . 
Ännu fler saknas . 
Överlevarna måste skyddas . 
Gilmore , hur snart kan du använda osynlighetsformeln ? 
Det finns inget kvar att dölja . 
Drakarna vet att vi är här . 
Du har den där blicken . 
Vad är det , Percival ? 
Ripley kände till var Whitestone låg hela tiden , men valde att säga det nu till Thordak . 
Jag tror jag vet varför . 
- Återstoden . 
- Hela Whitestones lager är stulet . 
Hon använde attacken som täckmantel när hon plundrade våra lager . 
Ripley har sinne för maskiner , inte magi . 
Vad ska hon med återstod till ? 
Jag har en teori . 
Thordak känner till platsen nu och Raishan vet att den är oskyddad . 
Om vi ska få tag i Ripley , måste det ske snart . 
Scanlan kanske kan hitta henne med mytsnidaren ... Om han var här . 
Jag kan kolla med mina kontakter i skrået . 
Om någon vet hur man fångar en orm så är det tjuvskrået . 
Behövs inte . Jag har henne . 
Obsidiantermit , en sällsynt sten svedd av gudomlig eld under katastrofen . 
Den kan bara hittas på en plats , Glintshoreön . 
Hon lämnade den medvetet . - En inbjudan . 
- Ja . 
- Men vi åker dit ändå . 
- Jag ser inget problem med planen . 
Älskling , jag vet att det är personligt för dig . 
Är du säker att du kan lägga band på dig ? 
Du sa att jag är förändrad . 
Låt oss hoppas på det . 
Vi ger oss av i gryningen . 
Okej . På tal om annat , var är Scanlan ? 
Han har förhoppningsvis mer tur än vi . 
Kaylie ? 
För sent . 
Du låg inte i sängen i morse . 
Jag fick smyga ut innan någon vaknade . 
Det har varit trevligt att ha något som bara är vårat , men det kommer en tid då man inser vad som är viktigt . 
Vill du berätta för dem ? 
Jag vill att vi är ärliga med varandra . 
Det vill jag med . Men att berätta kommer att förändra saker . Och de behöver vara fokuserade på uppgiften . 
- Du har nog rätt . 
- Självklart . Jag har alltid rätt . 
Titta på dem . Beter sig som om vi inte vet . 
Eller hur ? Hur dumma tror de att vi är ? 
De besudlade alla rum i Scanlans slott . 
Jag hörde dem stötande på biljardbordet ... Vi fattar . 
Trinket , du får stanna här och vaka över Cassandra och Whitestone . 
De behöver dig , förstår du ? 
Okej , vi känner inte till ett träd i Glintshore . Och Allura kan inte teleportera oss för vi kan hamna i havet . 
Så båt då ? 
Nej . Vi flyger . 
Resa ! 
Vill du ha min rock ? 
Tack , älskling . Men jag tror att vi är framme . 
Tack och lov . 
En hel dag utan öl . 
Jag är utsvulten . 
Oroa dig inte . Det finns nog en taverna runt nästa uråldriga , förstörda krök . 
Jag ska förstöra din uråldriga krök . 
Vänta här . Percy och jag sonderar terrängen . 
Jag ser inte ett skit . 
Tänk om det blir bättre ? 
- Vad ? 
- Om vi berättar om oss . 
Inte troligt . 
Scanlan kommer att reta mig obevekligen . 
Keyleth lär kalla mig hycklare . Min bror , jag kan inte tänka mig vad han skulle göra mot dig . 
Är det verkligen därför du är emot det ? 
För att skydda mig ? 
Varför är det så viktigt ? 
Behåll den tanken . 
Vad är det ? 
Vi berättar för de andra . 
Luftvägen är för riskabel . 
Ja . Men om det är någon där ute , så ser vi dem inte . 
Om det är någon där ute , så ser de inte oss . 
En stig . 
Så smidigt . 
Och säkert full av fällor . 
Jag lånar den lite . 
Varför spränger du inte din egen frukost ? 
Jag har en . 
Ett meddelande från Ripley . - De Rolo-vapnet . 
- Något är fel . 
Det var lätt . 
- Nästan ... 
- Nästan för lätt . 
Förlåt . Jag har alltid velat säga det . 
Det lät riktigt coolt . 
Vax är nästan klar . 
När vi når grottan , borde vi vara redo ... 
Det finns en anledning till att jag pressar dig om det här . 
Jag älskar dig . 
Percival , jag ... - Jag ... 
- Desarmerad . 
Kom igen , vi går . 
Stubby , kom igen . 
- Det är tyst . Nästan för ... 
- Nästan för tyst . Förlåt . 
Såg ni någon när du och Percy sonderade ? Vex ? 
Nej . 
Ja , menar jag . 
Ja , det var några vakter , de såg ut som sjömän . 
Percival . 
Orthax . 
Vax ? 
Vax ! 
Mor ? 
Vem gjorde det här ? 
Du , Vex ' ahlia . 
Din kärlek dödar . 
Percy . 
Fan ! 
Hallå , Percival . 
Du är sen . 
Välkommen till din fabrik . 
En produktion som drivs av ett magnifikt batteri som kombinerar det hemliga med Kabalens död , ånglokomotiv och Whitestoneåterstod . 
Allt inspirerat av din design . 
Så det är det du har sysslat med , utöver att förstöra mitt hem . 
Jag gjorde dig en tjänst . 
Du har alltid avskytt dina adliga plikter . 
Hur vågar du ... Och när min förvirringsgas tar sig in i dina vänners sinnen , är du fri från förpliktelser . 
En nystart för vårt partnerskap . 
Efter Whitestone är du galen om du tror att jag vill ha med dig att göra . 
En mindre olägenhet . 
Jag fick improvisera när jag insåg att skölden var falsk . 
Enda problemet är kraftkällan , en gång i timmen , som ett urverk . 
Se på dig . 
Försöker redan lösa det . 
Varför kämpar du emot , Percy ? 
Spänningen med upptäckter , ambitionen , det här är den du är . 
Jag har förändrats . Jag har blivit av med Orthax . 
Ett kostsamt misstag för dig . 
Men det här partnerskapet är obrytbart . 
När vi hittade varandra gjorde jag inte motstånd som du . 
Jag välkomnade insikten , klarheten , makten . 
Jag accepterade den jag är . Och jag är mycket starkare för det . 
Orthax kommer att få själarna av de som dräpts med dina vapen . 
Och i gengäld får alla egen makt . Och det blir upp till dem hur de nyttjar den . 
Men till vilket pris ? 
Din själ ? 
Magikerna tog båda våra familjer . 
Det var inte hämndlystnaden som drog Orthax till oss , det var därför vi drogs till Orthax . 
Du har rätt . 
Jag har lurat mig själv . Insisterat att jag har gått vidare . 
Det kanske är dags att acceptera att vissa sår inte läker . 
Jag känner till det allt för väl . 
Det gör vi båda . 
Vi är väldigt lika , Anna . 
Jag är inte perfekt . 
Men mina brister gör mig inte svagare . 
De gör mig till den jag är . 
Gå ! Ta honom ! 
Jag sa ju att han var värdelös . 
Låt mig ta hans själ . - Okej . 
Det är dags att avsluta vårt avtal . - Dags att avsluta vårt avtal . 
Sluta ! 
Evigt ljus ? 
Jag varnade , hon är inte där . 
Gudarna lovade guld och gröna skogar , att vara vid din sida . 
De ljög . 
Släpp mig . Släpp ! 
Vill du hjälpa dina allierade ? Frigöra dem ? Vill du det ? 
Tro i så fall inte på någon annan än dig själv . 
Sanningen finns i ditt blod . 
Kiki ! 
Fan . 
Vax får det att se så lätt ut . 
Det här tjänar ingenting till . 
Våra vapen är redo att skickas ut . 
Jag avslutar det du inte kunde . 
Vi skulle ha alla oskyldiga livs blod på våra händer . 
Jag tänker inte vara medskyldig . 
Framstegen kan inte stoppas . 
Snälla . Lämna mig inte här . 
Snälla ... Döda ! Alla är döda ! 
Va ? 
Fungerade det inte ? 
Pike ? 
Tack . 
Nej . Mor . 
Snälla . 
Jag hörde skrik . 
Mor . 
Jag kan behöva hjälp med den store . 
Ett bibliotek ? Ord ? Bara ord ? 
Varför finns det inga bilder ? 
- Pikey . Skadade jag dig igen ? 
- Nej , kompis . 
Jag är bara helt jävla slut . 
Vänta . 
Var är Percy ? 
Gömmer vi oss som en fegis ? 
Dina vänner är inte här och räddar dig , Percival . 
Svartkrut ? 
Ingen bra plats , de Rolo . 
Du har haft många chanser att döda mig . 
Svaghet kommer att döda dig . 
Sju ... 
Percival ! 
Vänta , Orthax ! 
Alltid smart , Percival . 
Och nu är hämnden din . 
Du kan se mig brinna . 
Jag är klar med hämnd , Anna . 
Dina överträdelser har förstört många liv bortom mitt . 
Vi förtjänar rättvisa . 
Jag förstår inte . 
Varför visar du nåd ? 
Jag vet hur demonen känns . 
Hatet som bränner i ådrorna . 
Jag kan hjälpa dig bli av med Orthax . 
Efter tid och botgöring kan du hitta en bättre väg . 
Din hjärna kan bli en gåva till världen . 
Du menar allvar . 
Vex . 
Percy ! 
Så upptagna Vilket håll skulle de gå åt Bandet mellan dem kändes evigt 
Skulle kärleken vinna Om de kunde ta det lugnt 
Med förvridna hjärtan och faror ... Nej ! 
Men livet går fort Och något kändes fel Hon sprang till honom Men han var borta 
Nej ! Pike ! 
Låt honom andas igen Han är borta . 
För nu finns inget kvar Vi kanske aldrig blir desamma 
Det var inte så det skulle sluta Snälla lämna mig inte . 
