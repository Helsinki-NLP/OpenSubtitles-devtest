Hon är en stråtrövare . Hon sägs vara beväpnad och extremt farlig . 
Vad har du gjort för att förtjäna en sån belöning ? 
- Hon dödade honom ! - Nej . Det var han ! 
Efter henne ! 
Jackson måste dö . 
Ödet har fört oss samman , Sofia . 
Dina förmågor har förbättrats . 
Jag är redo att lära mig mer . 
Bry dig inte om honom . Han är farligt . Giftigt . Drottningen är en förrädare . 
Du är jakobit . 
Halva Annes riksråd håller med mig . 
Isambard Tulley greps i Slough . 
Inser du att du hängs om jag inte ordnar det ? 
Det är vårt fel , så jag ska frita honom . 
Vi skickades hit för de här stackarnas skull . 
Är du verkligen Nelly Jackson ? 
- Åh , Nelly ! - Ut , allihop ! 
Tråkiga jordbor . Värsta förvirringen . 
Du kommer att dö , Nelly Jackson . 
Sofia ? 
Jag gillade din pjäs . 
Välsigne dig . Var är den andra ? 
Det här är en berättelse om passion och elände med en kvick hjältinna , Polly Honeycombe , som , inspirerad av hennes överlevnad efter ett brutalt rån , använde sig av den grubblande mr Scribble . 
Två som tillsammans trotsar sin hjärtlösa fars vrede , ignorerar hans önskan att förbjuda giftermålet och i enlighet med alla stora romanser kasta försiktighet , konventioner och anständighet åt sidan och rymmer . 
Jag måste erkänna att efter kärlekens första vågskvalp visade sig den ädle , eteriske mr Scribble vara mer hårig än väntat . 
God morgon , min kära . 
Kan det finnas stråtrövare här ? 
Inte en enda . 
Er vackra hjältinna fann att tankarna oåterkalleligt drev till ett ögonblick och en viss skurk med mycket mindre hår . 
Men med sin karakteristiska charm och optimism , försäkrade sig er hjältinna om att äventyret väntade . 
Men det visade sig snart att rymningar har vissa nackdelar , kära läsare . 
Som inte ett enda rån , städning utan en missförstådd bandit i sikte , och att upptäcka sin favoritklänning på en servitris . 
Min garderob är distinkt och jag skulle känna igen den överallt som den som stals av min stråtrövare . 
Åh , mr Scribble . Mitt rykte . 
- Vi är praktiskt taget gifta . 
Jag mår inte bra . 
Det var då en tanke slog er hjältinna som en blixt från klar himmel . 
Stråtrövaren som stal mina kläder gjorde det av kärlek . 
Det var så uppenbart . 
Tösen där nere är stråtrövarbrud . 
Genom att ge henne mina kläder , försökte han skapa en blek kopia av mig . Men ms Honeycombe kan inte ersättas . 
Jag fick förhöra henne . För mitt hjärta tillhör nu obestridligen min kärlekskranka stråtrövare . Och jag ska inte ge mig förrän ... Ack ! 
Er hjältinna svimmade - på ett tragiskt sätt när ... - Vänta . 
Du ska skriva ett lösenbrev , inte en jäkla roman . 
- Jag försöker ... - Kan vi ta tillbaka henne ? 
Vad säger vi till Japhia ? 
Att Amorous är en idiot . 
Jag är rädd att i en utsökt ironisk vändning , har skurkarna råkat kidnappa precis rätt person . För jag , miss Polly Honeycombe , är stråtrövarens sanna kärlek . 
Du menar väl inte vår Nell ? Nell Jackson ? 
En förkortning av Nelson , antar jag . 
Nell är ingen man . 
Hon är min syster . 
Det var därför de tog mig . 
De måste ha trott att du var Roxy . 
En stråtrövar ... kvinna . 
Är du helt säker ? 
Håll tyst om du vet ditt eget bästa . 
Skriv klart lappen . 
George här . 
Jag och " Polly Honeydrone " har kidnappats av luffare . De trodde att hon var du . 
Vi är i en lada utanför Uffington där de byter vår återkomst mot Nell . 
Pengarna eller livet . 
- Jag ? 
- Ja , du . 
Newgatefängelset hade ditt namn . 
Först Herne , sen det där . Något är på gång . 
- Som vad ? 
- Något mörkt . 
- En magiker kanske vill stoppa dig . 
- Varför ? 
De kanske gillar det hela , där sprättarna tror att de kan göra vad de vill mot vanligt folk . 
Det kan de inte . 
Det som pågick där är inte rätt . Vissa var mindre än George . - Det var fel . - Ja . 
Det behövde förändras . 
- Det kanske är därför jag har dig . 
- Ja . Jag ska nog inte till Amerika . 
Vi ska nog stanna här . 
Håller du med mig ? 
Nej . Vi ska inte rusa in i något . 
Vem som helst kan resa jorden runt och spränga folk , vi . 
Vi ska stå upp när något är fel och banka lite vett i dem som tjänar på misär och smärta . 
Ja . 
Ja . Okej . 
Okej . 
- George och Roxy då ? 
- De är säkrast i Abingdon . 
Är vi överens ? 
Vi ska rädda världen . 
Lugna nu . 
Vi börjar med kontinenten eller England , eller bara Tottenham . 
Jag trodde att ni var magiska . 
Varför kidnappar ni folk ? 
Vi var en riktig trupp . 
Vi var på Drury Lane , men ... Recensionerna var dåliga . Japhia förlorade sin roll . 
Och ? 
Så han slog halvt ihjäl ersättaren . 
Hela truppen smutskastades . Ingen ville ha oss efter det . 
Nu är vi häckkrabbor som knappt klarar sig och nu med ett barn på väg . 
Allt han vill är att bli känd , applåderad som han blev . 
De här showerna är flera år gamla . 
- God morgon ! 
God morgon . 
Lyd , så gör han er inte illa . 
God morgon , gamla pålitliga ... God morgon . God morgon . God morgon . 
Du ... Du har ... En bonde hade farhågor om att låna ut sin lada till vårt framträdande . Men vi har löst det nu . 
Varför har den stackars duvan fortfarande den här på sig ? 
Vi skulle ... Vem är det här ? 
Amorous . 
Amorous , din dumma idiot ! 
Vänta ! 
Hon hade klänningen . Hon hade den . 
Vilket muskedunder , va ? 
Nu har vi henne att göra oss av med . 
Min pappa är väldigt rik . 
Hur rik ? 
Han säljer peruker . 
Alla har peruker . 
Det är ju bra . 
Jag antar att vi inte ska döda dig än . 
Bäst att hon inte är sen . 
- Kom igen . 
- Farbror Jack ! Farbror ... 
Vi stöttar dig , Nell . 
Han ska hämta hjälp åt George . 
Varför ? Vad är fel ? 
Hon blev bortförd . 
Jag är så ledsen , Nelly . 
Vad menar du med bortförd ? 
- Nell ? 
- Har nån tagit George ? 
Några luffare . De vill ha dig , Nell , i utbyte . 
Sprätten läste lösenbrevet . 
De har även hans trolovade . Ja . Det är bäst att jag går . 
- Älskar du henne ? - Ja . Självklart . 
Kärlek och omständigheter hänger inte alltid ihop . 
Fegis ! 
Vi måste gå , Nell . 
De har haft George hela natten . Farbror Jack hittar inte hjälp i tid . 
Vi kan åka direkt till Uffington . 
- Jag behöver en häst . - Becky , häst . 
- Och till mig . 
- Nej . - Jag kommer . - Nej ! 
- Var är Rasselas ? 
- Vet inte . Vilket håll ? 
Nell ! - Vad gör du ? 
Gå tillbaka ! 
- Jag hjälper ! 
Va ? Nej ! Gå tillbaka , Roxy ! 
Sakta ner ! 
Vänta , Nell . 
Jag kan inte . Värdshuset är inte säkert . 
Det här är inte säkert . 
- Var är Rasselas ? - Han stack . 
Det gjorde han inte . 
Roxy , det var ... Det var ett upplopp och en stor mur kom emellan oss . 
Jag svimmade . 
Jag letade efter honom , men London är enormt , Roxy . 
Men när vi är åtskilda rasar allt samman . 
Nu hämtar vi George . 
- Vi är bättre tillsammans . Okej ? - Okej . 
Godolphin . 
Poynton ! Du har återhämtat dig . 
Hennes Majestät har saknat er frånvaro . 
Hon behöver lojala män . 
Jakobiterna kommer att dra nytta av Newgate . Allt detta kaos . Det har alltid slagit mig hur mycket du föraktar dem . 
Jakobiterna är giriga hycklare . 
De vill regera genom en marionett på tronen . 
Ett barn , en främling i England . 
Och de finns ibland oss , Poynton . Till och med i kronrådet . 
Berätta om du hör nåt . 
Självklart . 
Jag hörde talas om en förrädare . 
En som skickar brev till Frankrike . 
- Vem ? 
- Det vet du nog . 
Lord Godolphin , Poynton ... 
Vad ska det här betyda ? 
Är det sant ? 
I hans skrivbord . 
Inte mitt väl ? Det är ett misstag . 
- Berätta ! 
- Jag hoppades att jag hade fel . 
Poynton ? 
- Vad ? - Kom igen . - Släpp mig ! - Flytta på dig . 
The Courant borde göra fler intervjuer . Bättre ! 
" Ganska artig ? " Intervjua mig . 
Hon kunde ha dödat mig . Jag såg hennes ansikte . 
Valerian , håll upp hans huvud . 
Skoningslösa varelse . 
- Jag kan ta med det i The Medley . - Ja . 
Valerian , stötta hans huvud . 
Weekly Journal kanske medger att hon hade en viss sjaskig elegans . 
Sätt fart . 
Det finns en risk att Nell Jackson går under jorden , och det duger inte . 
Landet är i kaos . 
Folk vill ha heta nyheter . 
Och hon är allt de vill läsa om . 
Så vi behöver något som får henne att stampa runt igen . 
Idéer ? 
" Jackson äter bebisar . " 
Det har gjorts . 
" Vårtspridare " ? Nej , Valerian . Vulgärt . Man måste balansera djärva och exceptionella modeval med subtilitet . 
Annars , vad är man , förutom tafatt . 
Åh , nej . Nelly Jackson bryr sig inte om det . 
Jag kan hennes typ . 
Ja . 
Det här . Det här kommer att få fart på henne . 
Vad gäller min trolovade ... The Courant får rapportera , att eftersom han är den enda fången som inte har rymt från Newgate , är det ett uttalande om hans oskuld . 
Medan The Medley undrar om han är för dum för att hitta ut . 
- Eularia ? - Ja ? 
Nej , jag vill inte ha dessert . 
Du vill nog höra det här . 
Försvinn , sa jag ! 
Varför satte du mig i detta rum ? 
Du är lord Blancheford nu . 
Du borde ha lämnat mig i London . 
Du var ensam när mina män hittade dig . 
Ska jag beskriva ditt tillstånd ? 
- Allt är bra . 
- Inte alls . 
Inget blir bra igen på grund av dig . 
Nej , Thomas , inte på grund av mig . 
Hade nån annan gjort det ? 
- Du manade på mig . 
- Och du gjorde det ! 
Insikten att vi kan få allt vi vill ha ... om vi är beredda att göra vad som helst för det ... 
Vissa ser det som obegränsade möjligheter . 
Medan andra bara ser ... Skräck . 
Nej , nej , nej . 
Gör det inte . 
Jag förstår . 
Det gör jag . 
Och jag är rädd att jag måste be om ursäkt , Thomas . 
Du står inte ut , va ? 
- Nej . - Okej . 
Tänk om jag sa till dig ... att jag kunde få det att sluta på ett ögonblick ? 
Skuld . Skam . 
Vet du vad de bottnar i ? 
Ansvar . 
Du kan släppa det . 
Ni kommer att märka , käraste gnagare , att det inte är klokt att ignorera Isambard Tulley . 
Och att vi alla har vårt pris . 
Så kan ni sluta avbryta mig ? 
Om ni bara ... Lady Eularia ... Vem pratar du med ? 
Änglarnas ängel . 
Jag försökte bara träna en charmig liten mus . 
Ingen har besökt mig . Nya kläder till rättegången ? 
Som Valerians lille vän säger har flyttats till i morgon , eftersom du på nåt sätt har lyckats bli den sista fången i Newgate . 
Strålande nyheter , frigiven i förtid . 
Du har ordnat allt . Du har smörat för alla som behöver smöras för . 
Den här tiden i morgon planerar vi bröllop . 
Eller så är du död . 
Din lilla vän har släppt lös kaos . 
Så makthavarna har utövat sin makt . 
Och om domen är skyldig hänger de dig omedelbart . 
Men pengar är fortfarande allt . 
Säg inte att domstolarna är lagliga nu . 
Jag måste gå . 
The Medley gör ett specialinslag om dina brott och det säljer snabbare än vi kan trycka det . 
Eularia ? 
Hej då , Charles . 
Earlen av Godolphin greps som jakobit . 
Godolphin ? 
Brev hittades bland hans saker . 
Han är kapten för drottningens livvakt . 
Precis . 
Och nu är han gäst i Towern . 
Hennes Majestät vill att jag besöker henne . 
Gardet överlämnas nog till mig . 
Tänker du använda dem ? 
Jag ser till drottningen , så att James trupper kan avancera fritt . 
Vad står det i tidningarna ? 
De hävdar att landet står på randen till revolt . Att fängelset invaderades av Nell Jacksons folkarmé . 
Oavsett om de vet att det var du , så skakades London . 
Mår du bättre ? 
Jag mår utmärkt . 
Visst är det underbart ? 
Berusande . 
Ja . 
Jag hade nästan Jackson . 
Det får du igen . 
Du jagade iväg henne . 
Besvärjelsen utvecklades . Fängelset tog över . 
Håret vi använde brann upp . 
Vi hittar henne . 
Jag undrar om du förstår hur begåvad du är , hur viktig . 
Sån makt är inte för Nell Jackson . 
Det finns sätt att hantera henne . 
Okej , jag är här . 
Välkomna , mina damer och herrar . 
Var är min syster ? 
Vi har en speciell överraskning i dag ! 
Den hemska , den onda , den blodtörstiga , den djävulska , Nelly Jackson ! 
Vad i ... ? Ni är här för att bevittna historia . Nelly Jacksons tillfångatagande och fall av den oförliknelige ... Den stilige , hjältemodige , magnifike , mästerlige , underbarnet , geniet , virtuosen ... Japhia ! 
För dagens speciella framträdande har en plan kokats ihop . 
Ett utbyte . Nell Jackson mot sin lillasyster . 
Var är hon då ? 
" Måste du bränna ut båda mina ögon med heta järn ? " 
" Jag måste . Måste . " 
Shakespeare . 
- Jag har läst mycket om dig . - Jaså ? 
Omöjlig att besegra , sägs det . 
Omöjlig att skada . 
Men det är hon inte . 
George . 
Stå still . 
Vi skulle inte skada henne . 
Lägg ner den , jag gör som du vill . 
Ni lyckostar ska inte bara få bevittna gripandet , utan även avrättningen av ett av vår tids monster . 
Anklagelserna stämmer inte . 
- Jag är inte ... 
- Det är oväsentligt . Det är vad du uppfattas som . 
Dödar jag dig är jag en hjälte . 
Jacksons bägare innehåller gift . 
Vi skålar för hennes frånfälle . 
Det spelar ingen roll hur stark eller snabb demonen inom dig är , Nelly Jackson . Jag tvivlar på att den kan rädda dig från odört som du dricker själv ! 
Det är den andra . 
Det är lugnt , va ? Om jag dricker ? 
Vi testar inte . Jag ... 
- Vad ? - Jag vet inte , Nelly . Jag är bara människa . 
Gör nåt då . 
Distrahera honom . 
Gift ? 
Den gamla godingen ? 
- Bu ! - Det är en klassiker . 
De kommer att berätta vad du har gjort och du hamnar i snaran . 
Det beror på vinkeln , eller hur ? 
- Tidningarna gillar inte dig . 
- Jag är oskyldig . 
Jag är trött på att se dig i varje tidning . 
Ditt ansikte där mitt borde vara . 
Du kommer att vara död och jag känd . 
Släck lampan ! 
Kära nån . 
Den stora Japhia ser svettig ut . 
Tycker ni inte det ? 
Stick ut ett av den lilles ögon . 
Stick ut båda två . 
De funkar ändå inte . 
Okej . 
För ödet . 
Ja . Skål . 
Hej då , Nelly Jackson . 
Nej , nej , nej . Nelly , nej . 
Nej , kan inte ... 
Klantade jag mig ? 
Jag svalde en fluga . 
Är du okej ? 
Bara bra . 
Döda dem ! 
Mina sista ord . 
- Vi behövde inte höra dem . - Bra gjort . 
Det var det bästa jag har sett på åratal . 
Lycka till med det . 
Kom igen . Nu går vi , Roxy . 
En av militärfruarna fick barn under en marsch . 
Hon gick till vägkanten och klämde ut det bakom en buske . 
Jag säger bara det . 
- Det var omtänksamt . 
Och det snöade . 
Hon hann ikapp oss vid lunchtid . 
Väldigt anständigt . Inget strul . 
Födelsens mirakel är inget för mig . 
Vad tycker du om titeln " Rebelliska Nelly " ? 
Jag hjälper dig inte skriva en pjäs om mig . 
Det finns nog med strunt . 
Jag vill att du ska veta , att det kvittar att din far var tjuvskytt . 
Det var han inte . 
Visst . Självklart . 
- Vad står det mer ? Vad mer ? - Inget . 
Nej . Vad ? Berätta . 
Uppenbarligen förtal . Uppenbarligen . 
Weekly Journal Nell Jacksons slyngelfamilj . Men de säger bara , att äpplet inte faller långt från trädet . 
Hela familjen är rutten . Att de också är tjuvar och i allmänhet inte bättre än de borde vara . 
- Jaså . - Du vet hur de skriver om kvinnor ibland . 
Det kvittar . 
Folk tror inte på det . 
Nej , det är precis vad folk kommer att tro . 
Okej . 
Vi ska slå sönder pressarna . 
De bygger bara fler . 
Ingen kanske har trotsat dem förut . 
De där blaskorna livnär sig på elände och gör det värre . 
De skapar monster som snigeln Japhia och ljuger . 
Vi måste visa att de inte kommer undan . 
Folk måste få veta att sanningen spelar roll . 
För det gör den . 
Vi kan stoppa dem . 
Det är nog meningen . 
Ja . Okej . 
Okej . 
Kom igen . 
Kan vi leta efter mr Rasselas också ? 
Kan du skjutsa oss ? 
- Sofia . 
- Rasselas ? 
Jag har försökt nå dig . Jag måste prata med dig . 
Är hon här ? 
Nell ? 
Nej . 
Jag var på Newgate . 
Var du ? 
Hur var det ? 
Jag läste om det i tidningen . 
- Blev du skadad ? - Jag tyckte ... Vad ? 
Att jag hörde din röst . 
Vad sa jag ? 
- Hur lät jag ? - Jag vill veta varför , Sofia . Och den där killen är här . 
Greven av Poynton . 
Han sitter i riksrådet . 
De rör sig i såna kretsar . De är annorlunda . 
Kanske för dig . 
Vad gör han där ? 
Han är en vän . 
Har han en hållhake på dig ? Du kan berätta för mig . 
Han har bara hjälpt mig . 
Och jag har alltid kontroll . 
Jag hade nog med kontroll i Newgate . 
Valde du att göra det ? 
Det var monstruöst . 
Det var monstruöst att överge mig när jag behövde dig som mest . 
Natten då min far dog , kastade du bort all vår historia . - Vilken historia ? 
- Vilken historia hade vi ? 
- Du är min vän . 
Sofia , din far köpte mig ! 
När du blev för gammal , skickades jag till stallet som en gammal leksak ! 
Jag behandlade dig aldrig så ! 
Du var vänlig och stod mellan mig och Thomas . Jag är tacksam . Men det var aldrig ... Jag var aldrig här frivilligt . 
Du kan få slut på allt det här . Säg bara sanningen . 
Vet du inte vad de gör med Thomas om de får reda på det ? 
Han är min familj . 
Nell , då ? Hennes familj ? 
Minns du när Thomas brukade fånga grodyngel , skalbaggar och spindlar ? 
Och du och jag släppte dem fria . Om han försökte straffa mig , stoppade du honom . 
För du är rättvis , Sofia . 
Gå till henne . 
Gå tillbaka . 
Vänta . 
Du kommer att få sårröta . 
Lycka till . 
