Stopp ! Vad gör ... Hallå ! 
Okej . Dörren är öppen . 
Vilken av fångarna är det ? 
Jag sa ju det . Sektledaren . 
Stor belöning om vi får ut honom . 
Du där . Råkar du vara en sekterist ? 
Ursäkta ? 
De andra cellerna är tomma . 
Det här måste vara vår jävel . 
Letar ni efter den tokiga mystikern , missade ni honom med två dagar . 
Fångenskap gick inte ihop med hans konstitution . 
Ja . Äckligt . 
Fan . 
Där missade vi den belöningen . 
Kanske inte . 
Du verkar inte höra hemma på ett sånt här ställe . Lustigt . Det gör ni . 
Vi har lite ont om pengar och du pratar som om du är rik . 
Hur mycket skulle du vara värd ? 
En smärre förmögenhet . 
Om jag inte var pank för tillfället . 
En detalj du kunde ha undanhållit tills du var fri . 
Varför ljuga ? 
Ni upptäcker snart att jag är fattig . 
Jag är helt ensam i världen . 
Ni kanske kan relatera . 
När man når botten är sanningen det enda man kan köpslå med . 
Att erkänna att man behöver hjälp förändrar folks sympati . 
Du är kass på att förhandla , det vet du , va ? 
Men du är brutalt ärlig . 
Ni kan behöva den ärligheten en dag . 
Okej . 
Vi ser vart ärligheten tar oss . 
Vad heter du ? 
Whitestones befolkning är vana vid förlust . 
Sorg har blivit vår mest bekanta granne . 
Trots det är sorgen av den här tragedin grymmare än resten , då vår älskade bror , vän och nobla son har tagits ifrån oss på nytt . 
Likt hans familj , var Percival de Rolo en man med djup hängivenhet till sitt hem och lojalitet till sitt folk . 
Han var inte religiös , men han trodde på Whitestone med hela sin själ . 
Hans hjärta fann mening i vår historia , men hans sinne lyste upp vår framtid . Han ägnade timmar av sitt liv åt att snida vårt arv med tidens orubbliga stämjärn . 
När vi böjde oss stod Percy stark och påminde oss om att hoppet är en låga värd att vårda . 
Och trots att vi tar farväl idag , kommer Gryningsfadern att hålla hans låga vid liv inom oss alla . 
Vi ber i hans namn , för in ljuset där mörkret bor . 
För in ljuset där mörkret bor . 
Vad hände ? 
Var är Percy ? 
Det finns en anledning till att jag pressar dig om det här . 
Jag älskar dig . 
- Syster . 
- Jag kunde inte säga det . 
Jag var inte stark nog . 
Du är den starkaste jag känner . 
Jag var orolig för hur han och du skulle reagera . 
Jag stängde hjärtat när jag skulle ha öppnat det . 
Jag för otur med mig . 
Varför säger du det ? 
Min kärlek förstör allt jag rör vid . 
Tanken på att känna så starkt igen gjorde mig livrädd . 
Och nu får Percy aldrig veta . 
Såklart han visste . 
Han må ha varit en reserverad , retfull skit , men han var skarpare än mig . 
Och varje gång du såg på honom visste jag . 
- Gjorde du ? 
- Bara en dummer hade missat det . 
Och han var inte dum . 
Men det som blev osagt förblir det . 
Hur kan jag leva med det ? Hur kan någon det ? 
- Hej . 
- Hej . 
Är Vex okej ? 
Är du det ? 
Förlåt att jag stack . Från oss . 
Kom in . 
Framtiden har skrämt mig så länge . 
Men det är en framtid som ännu inte har skrivits . 
Och jag börjar tro att ödet blir vad man gör det till . 
Det är okej att vara rädd . 
Men vi kan möta allt , om vi är tillsammans . 
Jag vill inte vara ensam . Vill du ? 
Jag har inte heller velat vara själv . 
Det är inte ditt fel , Scanlan . 
Jag hade kunnat stoppa dig från att gå . 
Varför gjorde du inte det ? 
När alla alternativ är dåliga , följer man hjärtat . 
Jaså ? 
Vad händer om det misslyckas också ? 
Det finns fortfarande ett sätt . 
Vad fan vill du ? 
Beklaga sorgen . Och planera vårt nästa drag mot Thordak . 
Hur fan vågar du ? 
Vi har inget avtal längre , minns du ? 
En handfull av hans avkomma har redan kläckts . 
Dussintals följer inom kort . 
Om du inte vill att Tal ' Dorei förgås så som din vän gjorde , föreslår jag att vi återupptar avtalet . 
Vi behöver tid , vi sörjer . 
Min syster är en spillra . 
Jag ville inte betunga dig med det här , men det är dags att du får veta sanningen om din familj och Thordak . 
Vex , vi måste prata . Du ... Vad är allt det här ? 
Jag är oanvändbar för er just nu . 
Distraherad . 
Jag måste rensa skallen . 
- Trinket och jag campar ... 
- Vex ' ahlia , du kan inte . 
Smärtan du känner , det är inte första gången vi känner den . 
Va ? Vad säger ... Berättelserna om förstörelse som Thordak drar . Skrytet om städerna han brände . 
Hamnstaden Callavon . Gremedash . Byroden . 
Ja , er hemstad , om jag minns rätt . 
Mor . 
Ert öde har varit tjudrat till Cinderkungen sen ni var barn . 
Det är dags att ni slutar ignorera det . 
Thordak är ert öde . 
Den sorgen lamslog oss båda i flera år . 
Kanske hela våra liv . 
Och förlusten av Percy kan göra samma sak om vi tillåter det . 
Vad är det du säger ? 
Stubby , vi kan hämnas dem båda . 
Ett dussin omogna drakar förstörde Whitestone . 
Och enligt Raishan kommer Thordaks ägg snart att kläckas . 
- Om de gör det ... 
- Då är vi helt körda . 
Det skulle vara dåligt , ja . 
Jag litar minst på henne , men vi lyssnade inte på henne sist , och Percy dog . 
Men att ta Emon från världens farligaste drake . 
Ni har försökt förut . 
Om ni inte har gömt undan en armé , vad är annorlunda nu ? 
Tänk om vi hade en armé ? 
Jösses . Grog , jag sa till dig att inte äta Percys verkstadspasta . 
Nej , vi har fått vänner var vi än har varit . 
- Ja . Och fiender . 
- Jo , visst . Men om Thordak vinner kommer både vänner och fiender få lida . 
Det är större än Whitestone , till och med Tal ' Dorei . 
Han har rätt . 
Jag kanske kan övertala ashari om hjälp . 
Vi kan fråga Zahra och Kash i Vasselheim . 
Och Jordbrytaren Groon . 
Han är grym . 
En tilltalande idé , Grog . 
Men du pratar om några få krigare . 
Det räcker knappast . 
Vad sägs om tusen Syngornsoldater ? 
Det skulle göra skillnad . 
Vad väntar vi på då ? 
Fan ! Varför måste jag alltid vara betet , Z ? 
För , älskade Kash , du är så jäkla attraktiv . 
Det är helt rätt . 
Okej , vi släpar tillbaka honom för belöningen . 
Hur mycket kommer skrået betala för honom ? 
Hundra guld ? 
50 ? 
Nej . 25 . 
Vad sägs om att uppgradera till något fjälligare ? 
- Pratar du om drakar ? 
- Nej , nej . Nej ! Sist vi hjälpte er dog vi nästan . 
Kom igen , vill ni inte få upprättelse ? 
Eller åtminstone en större belöning ? 
Okej . Vi vet att vi står i skuld till er , men nära döden och en säker död är inte samma sak . 
Ursäkta . Jag och Z ? Paketavtal . 
På tal om det , var är din syster ? 
Så du lyckades . Fick tag i Fenthras båge . 
Har du kommit för att få mitt beröm ? 
Trevligt att träffa dig med , far . 
Men nej , jag behöver inte ditt godkännande . Jag söker något som är svårare att ge . 
Våra arméer ? 
Jag har hört att ni samlar styrkor , men jag är rädd att det är omöjligt . 
Thordak kan få Emon , för min del . 
Våra styrkor måste stanna här för att skydda Syngorn . 
Din militär är den enkla delen . 
Vad vill du då ? 
Jag vill att du erkänner sanningen . 
Draken dödade mor . Elaina . 
Jag har i alla år trott att hennes död var mitt fel . 
Att vi var skälet till att hon skickades till Byroden , och om vi inte hade fötts , hade hon kanske levt . 
Och vet du varför jag trodde det ? 
För att du trodde det med . 
Du beskyllde oss för hennes död . Struntprat ! 
Det har jag aldrig sagt . 
Du vände ryggen åt dina barn ! 
Du stängde ute oss när vi behövde dig . 
Vi fick klara oss själva i en värld som förtär kärlek och hopp . 
Det enda rådet du nånsin gav oss var att vakta våra hjärtan . Att inte släppa in någon . 
Och nu vet jag varför . 
Du var för stolt för att erkänna att du älskade henne . 
Hennes död sårade dig lika mycket som oss . 
Det är din sanning . 
Det var längesen . 
- Jag har gått vidare . 
- Inte jag . 
Du lärde mig att min kärlek var giftig . 
Jag lärde mig läxan så väl att jag höll en bra man som öppnade sig för mig på avstånd tills det var för sent . 
Och nu skulle jag ge allt för att få hålla honom , berätta vad jag känner , och att inte vara den känslokalla idiot som du skapade . 
Men allas smärta är deras egen . 
Och han är borta . 
Vex ' ahlia ... Förlåt . 
Det är det enda jag kan köpslå med , far . 
Sanningen . 
Om du har någon kärlek kvar för mig , eller mor , marschera då till Emon och bevisa det . 
Och om inte för oss , tänk då på dem som ska bo i den här världen när du är borta om det finns något kvar . 
Kash och Zahra nekade vår inbjudan . 
Räcker det här ? 
Jag är här . 
Vi möter det tillsammans , vad som än händer . 
Inte mitt öde . Inte ditt . 
Vårt . 
Vad gör du ? 
Att sjunga lugnar ibland mina nerver . 
" Kaylies sång . " 
Din text är jättefin , Scanlan . 
Har du visat henne den ? Nej . 
Och jag ska inte det . 
Jag försökte vara pappa och delaktig i gruppen och jag misslyckades med båda . 
Det kanske finns en lösning . 
Ja , det gör det . 
Inga fler distraktioner . 
Hörni ? Ni måste se det här . 
Kompaniet , stanna ! 
Herrejävlar ! Hon lyckades ! 
Framåt marsch ! 
Må han släcka lågan av hämnd och krig . Rulla tillbaka den ! 
Släpp ! 
Våra soldater är redo . 
Vad är attackplanen ? 
Vi ska driva ett tvådelat anfall . 
Din Syngornarmé , Groons krigare , och Whitestones vakter kommer att marschera genom stadsporten och ta sig an Thordaks avkomma . 
Med eldtämjare och luftashari framför för att skydda mot eldattacker . 
Allura och jag hjälper till med vår magi . 
Och medan markstyrkan tar sig an Thordaks avkomma , använder Vox Machina distraktionen för att nå hans lya . 
Hur tar ni er in ? 
Jag har sonderat . 
Vi tar oss in från luften . 
Det går inte . 
Hans barn vaktar den nu . 
Och vem är du ? 
Hon ... Jo ... En informant . Hon heter Larkin . Det är ett kodnamn . 
Det finns en oskyddad bakingång till Thordaks lya . 
En tunnel vid klipporna som är för liten för en drake . Men stor nog att ta sig in i . 
Och du försäkrar att tunneln är öppen ? 
Jag ger er mitt ord . 
Så vi dödar de små medan ni använder relikerna mot Thordak . 
Plus skölden . Om jag får den att fungera . 
Det ... Det är en bra plan , lady Vex ' ahlia . 
Men fungerar den ? 
Det måste den . 
Infanteriet , formera er ! 
Lycka till därute . 
Det är en ära att ha er på vår sida . 
Stormlorden är på er sida . 
Det är allt ni behöver . 
Är allt klart , Grog ? 
Vex , förlåt att jag inte var där . 
Jag vet , Scanlan . 
Efter idag kanske alla kan förlåta varandra . 
Är du redo , syster ? 
För Percy . För mor . 
För Exandria ! 
Fan . Ner ! 
Vi tar oss inte in där . 
Rök men ingen eld . Hur fungerar det ? 
Och inget motstånd . 
De borde ha upptäckt oss nu . 
Åtminstone mig . 
Vi har som tur är Raishans ingång . 
Om den inte är där ? 
Jag ser den . 
Landa där . 
Det är så mycket rök . 
Vi ser ingenting . 
Stanna ! 
Ynglingar ! 
Magiker till fronten ! 
Inta positioner ! 
Förbered ballisterna ! 
Varför attackerar de inte ? 
Känner ni det ? 
Helvete . 
Nej . Hon avslöjade oss ! 
Är den förseglad ? 
Den är varm än . 
Thordak måste ha smält den för cirka en timme sen . 
Grog , kan du slå igenom den ? 
Det kommer att låta en del . 
Jäklar . Jag är starkare än jag trodde . 
Det är nog inte du , grabben . 
Helvete ! Jag sa ju att vi inte kunde lita på henne . 
Vänta . Då betyder det ... 
Har han lämnat lyan ? 
Herregud ! 
Vad har jag gjort ? 
