Det har gått 500 år ... och Lautrecs skatt är fortfarande Neapels största olösta mysterium . 
Den ligger nergrävd djupt i stadens inre , och ingen har ännu lyckats att hitta den . 
Här är lagfarten för fastigheten . 
Lägenheterna står tomma om tre dagar . 
Sakta i backarna ... 
Var är den ? 
Kom igen ! 
Spring efter honom ! 
Nej , inte ni . Portföljen ! Hämta portföljen ! 
- Nu tar vi honom ! - Kom igen ! 
Vart tog han vägen ? 
Följ mig ! 
Du hoppar från tak till tak Folket skriker därnere Munaciello är tillbaka ! 
Stanna , din fähund ! 
Kom hit och ta mig . 
Killen är död . 
Vi sticker . 
- Sasà , rita honom utan hår . 
- Nej . 
- Sasà , han är skallig ! 
- Nej , sa jag ! 
Han hade krulligt hår senast någon såg honom . 
Stämmer inte det ? 
- Jag sa att han är skallig ! 
- Allvarligt ? 
Sluta nu ! Kom , Gennà , vi går hem . Mamma väntar på oss . 
Vi har bara några dagar kvar ihop . Vi måste ta vara på tiden . 
Sasà , man stavar " Wonderboi " med W. 
Det är så man uttalar det . Jag skriver som det låter . 
Det är en jaguar på skateboarden . 
Ska du börja nu också ? 
Wonderboy är inte brasiliansk som du . 
- Sluta . 
- Vad säger du ? 
Hörni , akta er ! 
- Aniè , vart ska din pappa nånstans ? 
- Ingen aning ... 
Kom . Vi gör klart teckningen sen . 
När då ? 
Har ni glömt att vi måste göra ritualen ? 
Kom igen . 
- Ja , nu går vi . - Kom . 
- Okej . Hej då . 
- Hej då ! 
Hej då . Vi ses . 
Ta den här , Terè . Annars mördar mamma mig . 
Kom nu . 
Vänta på mig ! 
- Har ni packat alla era saker ? - Ja ! 
Jaha ... 
Du är så vacker , älskling . 
När du gifter dig ska jag sy nåt ännu finare åt dig . 
- Nu börjar du igen ! - Nej ! Stå still ! 
Jag har bara tråcklat . Stygnen går upp . 
Tänker du på mitt bröllop , inte på att vi ska flytta om tre dagar ? 
Det är just därför . 
Pappa , inget kommer att hända med sonen till butiksägaren . 
Jag åker hellre till Tyskland och bor hos mamma . 
- Du säger ju att du inte vill flytta . - Ja , det är så man säger . 
Jag ska berätta en hemlighet för er ! Ser ni alla fina slingor i mitt hår ? 
Ni tror kanske att det är shatush , men det är det inte . 
Det kallas " bala-layage " . Balayage ! 
- Vad vill du , Aniello ? 
- Jag vill låna pappas scooter . 
Fråga din pappa ! 
Avbröt du mig när jag filmade för det ? 
Det som gick så bra . 
Gå nu , hjärtat . Gå ! 
Vad ? 
Vad menar du ? Det är mitt rum , pappa . 
- Får jag låna din scooter ? 
- Den är trasig . 
- Raffaele och Gennaro åker imorgon . 
- Lycklig resa . 
Vad gör hyresvärden här ? 
Det är inget . 
Gå och lek nu . 
Fru Angè , oroa er inte . Jag fixar det . 
Ja , det hoppas jag . 
ANDARNAS SLOTT Gennà , historien som jag lade upp har redan 20 kommentarer . 
De är alla från desperata tjejer . 
Hör bara : " När du är inte där , är jag rädd att gå förbi ditt hus . " 
Vad säger du om det ? 
" Adress i Brescia ? " Hon vill ha min adress ! 
Snyggt ! Men ingen av dem har dykt upp här . 
Är ni inte klara än ? 
Rafè , Gennà , kan ni skynda er på ? 
Vad skönt att vi flyttar imorgon . 
Äntligen lämnar vi den här skitiga stan . Vår nyårsafton kommer att bli den bästa någonsin ! 
Brescia ger oss allt som Neapel inte kan . 
Ni får en bättre framtid och er pappa får ett stadigt jobb där . Och vi slipper äntligen vår hyresvärd . Hon har bestämt över oss och vår hyra . 
Håller du på med Neapels hemsökelser igen ? 
I Brescia finns det inget sånt . 
- Inte ? 
- Nej , du behöver inte den , Gennà . 
Vet du vad vi gör ? 
Vi slänger den . 
- Vad säger du ? - Kom ! 
Och så packar vi färdigt . Eller hur , mamma ? 
- Bra . Seså . - Vart ska vi ? 
- Följ mig ! 
- Gå nu . 
Kom ! Ta med dig boken . 
Jäkla ungar ... 
Jag har slitit så för att få stipendium . 
Jag vill läsa arkeologi . 
Jag vill studera i Neapel . Italien är bästa stället för arkeologer . 
Jag tänker inte vänta på att vår hyresvärd sparkar ut oss . 
Sasà , vart ska du ? 
Ni ska väl inte hitta på några dumheter ? 
Jag ska bara säga hej då . 
Jag ska prata med vår hyresvärd . 
- Jag klarar inte den tonen ... - Nej , morbror . 
Du sjunger inte rent . 
Försök sjunga själv . Du vet att jag inte vill sjunga efter att mamma försvann . 
Varför vill du inte åka med mig på kryssningen ? 
Du behöver inte sjunga . Du får hänga med mig och säga till när jag sjunger fel . 
Jag vill inte prata om det här . 
Jag vill stanna här . 
- Hyresvärden slänger ut oss om tre dagar . 
- Sluta , nu . 
Jag ska bo hos mina kusiner . Jag stannar i Neapel . 
Statyetten . 
Ta reda på statyetten . 
Gör det genast . 
Donna Angè , killen är död . Han hoppade ner i Neapels djupaste brunn och han landade pladask . 
Ni blev grundlurade , idioter . 
Ni såg honom inte , han kan klättra uppför väggen . 
Han är inte mänsklig . 
Folk säger att Neapel har fått en ny Munaciello . 
Snacka inte strunt ! 
Munaciello är död . 
Du är en idiot . Om du inte får tag på statyetten till mig , skär jag öronen av dig . 
Jag förstår . 
Sätt fart . 
Du ande , vars hjälp jag söker ... Jag ger dig mina örhängen jag fick inför min första nattvard . 
Nu är de dina . 
Hjälp mig . Du vet vad jag önskar mig . 
Jag vill se mamma igen . 
Nåväl , jag hoppas att du gillar örhängena . 
Jag måste gå . Jag ska ta farväl av mina vänner . 
Men imorgon kommer jag med en ny gåva , okej ? 
Ni anar inte vad jag fått höra ! Jag är på väg , men ... 
Åh , nej ! Attans ! 
Nu går vi . 
Ni anar inte vad jag fått höra . Jag är på väg , men ... 
Vi får vänta på honom därnere . 
Han vet var vi ska träffas . 
Knäppgöken är därborta . 
Var tysta . 
- Kom . - Vart ska ni ? 
- Vi tänkte bada . 
- Bada ? 
I december ? 
Ni tänkte gå till Andarnas slott , inte sant ? 
Det är Neapels farligaste plats . 
- Håll er borta därifrån ! 
- Spring ! 
Aniello är inte här än . 
Alla måste vara här . 
Hans telefon är avstängd . Han klarar sig ändå . 
Än sen ? Han är vår kompis . 
Terè , vi måste börja . 
Sätt igång , Gennà . 
I sirenens namn , hon som alltid har varit vår beskyddare , bildar vi nu en pakt som förbinder oss för evigt . 
Siren Parthenope , vi överlämnar härmed den bok som vi har författat under våra glädjefyllda år ihop . 
Ta varandras händer . 
Om exakt fem år , när vi alla är gamla nog , kommer vi att återvända hit . Vi ska utforska alla hemligheter som finns i vår kära stad , vars historia spänner över 5 000 år . 
Till oss och Neapels hemligheter ! 
- Alltid tillsammans ! - Alltid tillsammans ! 
Wonderboy ! 
Jag har bevis på att han finns i verkligheten ! 
Han stal hyresvärdens statyett . Hon är besatt av den . 
Hon beordrade pappa att hitta den ! 
Det var därför han hade bråttom i morse ! 
Han tog statyetten till underjorden ! 
- Varför ska vi bry oss om det ? 
- Varför ? 
Hyresvärden vill ha tillbaka statyetten ! Vi kan utpressa henne om vi hittar den ! 
Ni slipper flytta ! 
Era hem i utbyte mot statyetten ! 
- Ta det lugnt . 
Hur ska vi hitta den ? 
- Den är i underjorden ! 
Vi har ritat kartor i fem år . Inte sant , Gennà ? 
Jo , men de underjordiska gångarna är över 40 mil långa . Och vi har bara utforskat några kilometer . 
Hyresvärden kommer inte att ge efter för nån utpressning . 
Ja ... 
Har du inte märkt hur hon behandlar oss ? 
Hon hatar barn . 
Menar ni allvar ? 
Ni är mina enda vänner som bryr er om mig ! 
Varför backar ni nu ? 
Du , Aniè ... Gör inte det här svårare än det redan är . 
Okej . Gör som ni vill . Då gör jag det här själv . 
Jag går in genom Gaiola . 
- Nej . - Aniello , sluta . 
- Aniello ! - Vart ska du ? 
- Aniello ! - Aniello ! 
Herregud . - Aniello ! - Aniè ! 
- Aniè , sluta ! 
- Nedrans ungar ! 
Jag visste att ni var här ute och hittade på dumheter . 
Vi måste snart åka härifrån . 
- Kom nu . - Vänta . Först ... 
- Säg inget ! 
- Gå och packa ! 
Vad gör han ? 
Börjar du nu igen ? 
Hem med er ! Skynda på ! 
- Har du inte hört ... - Vad ? Inte ? Såg du antikhandlaren Enzo ? Han gick just upp . 
- Jaså ? - Ja . 
Överlämnandet igår ... 
- Det blev inte av ... - Det var illa . 
Ja . Vi får se hur det här går . 
Vad vill du ? 
Eftersom du inte gav mig statyetten , får du inga lägenheter . 
Hade du gjort en uppgörelse med tjuven ? 
Du är en sån idiot . 
Det är du som måste ha snackat med någon ! 
Jag ? 
Du är en riktig klant . 
- Vad säger du ? 
- Släng ut honom . 
Släpp mig . Vad gör ni ? Rör mig inte ! 
- Håll tyst ! 
- Ingen får lura mig ! 
En deal är en deal . 
Jag ska hitta statyetten , och du ska ge mig fastigheterna . 
Stick härifrån , din idiot . 
Det här är inte över . 
Vad händer med våra hem ? 
Vad vill du ? Vem är du ? 
Jag förbannad ! 
Det här är inte över ! 
Vi provar här , Sasà . 
Chihuahua , godmorgon . 
Vi letar efter Aniello . 
Vi behöver veta var han är . Det är nåt som har hänt . 
Ni anar inte vad som hänt mig . 
Men Aniello är inte här . 
Ni får gärna leta reda på honom . 
Stick och lek , nu . 
Kom igen ! 
Det är vi . Öppna . 
- Aniello är inte hemma . 
- Attans . 
Han tog sig ner under jord för att leta reda upp Wonderboy . 
Ska vi ringa polisen ? 
- Har du redan blivit nordbo ? 
- Vi måste prata med hans mamma ! 
De bryr sig inte om honom . 
Då går vi själva ! 
Är du galen ? 
Utan hjälp ? 
Kan vi inte be knäppgöken att hjälpa oss ? Clemente ! 
Han vet allt om stans undre historia . 
Han är också ganska knäpp . 
Sasà har rätt . Det är vår enda chans . 
Aniello slängde sig från klippan för vår skull . Vi ska rädda honom . 
- Raffaè ! Gennà ! 
- Följ mig . 
- Är ni klara med packningen ? 
- Ja , nästan ! 
Kom . 
Raffaè , vad är planen ? 
Packa era ryggsäckar . Vi ses på det vanliga stället . 
Vem är du ? 
Hur kom du hit ? 
Jag är vilse . Jag hoppade i vattnet och så kom jag hit ! 
- Var hoppade du i nånstans ? 
- Vid Andarnas slott . 
Kom du hit från Andarnas slott ? 
- Varför då ? 
- Tänker du inte hjälpa mig ? 
- Hjälp mig ! 
- Rör dig inte ! 
Vad gör du ? Vart tar du vägen ? 
Herregud . 
Så du är ... 
Du kan säga som det ligger till . 
Du är Neapels nya Munaciello . Du stjäl från rika och ger till fattiga ! 
- Ja , jag är Robin Hood . 
- Nej ! 
Du är bättre än Robin Hood . 
Du är Wonderboy . 
Jag heter Tonino . 
Vi har stängt . 
Så du är min nya hyresvärd ? 
Vad vill du mig ? - Följer du efter mig ? 
- Varför träffade du vår hyresvärd ? 
Varför ska du hitta hennes statyett ? Vad handlar det om ? 
Det är inget viktigt alls . 
En kille på skateboard körde förbi mig och stal den . 
- Vilken kille ? 
- Jag sa att vi har stängt . Ge dig av nu . 
Stick . 
Stick ! 
Etthundratjugoett trappsteg ... 
Ja , men vi såg så många fantastiska saker där nere . 
Ja . 
Och alla stegen är värda det här . 
- Eller hur , Maltè ? 
- Naturligtvis . De gör inget om det är 150 . 
Jag är väldigt nyfiken . 
Jag vill höra mer om historierna du berättade . 
Det är en fantastiskt värld därnere . 
- Vi har några böcker här som ni kan ... 
- Jag gillar inte att läsa . 
Vi har dvd-skivor också . 
- De gillar jag inte heller . 
- Hur kan jag hjälpa er ? 
Du ska själv berätta om stadens legender för mig . 
Släpp mig . Låt mig vara ! 
Bäste doktorn ... Nu ska du få berätta en trevlig saga för oss . 
Vad ? 
Jag är större än du . 
Hördu ! Låt mig få lite andrum . 
Jag måste fokusera på att hitta rätt . 
Hitta vägen ut , menar du ? 
Så här ligger det till : Jag vet inte hur jag hamnade här . 
Nu ska jag hitta en väg ut . Sedan går du din väg och jag min . 
Är det uppfattat ? 
Okej ? 
Jag är bara nyfiken ... Du har byggt om din skateboard , va ? 
Jag borde ha lämnat dig däruppe . 
- Hur lyckas du skaka av dig alla ? 
- Vad då " alla " ? 
Vad snackar du om ? Du är en superhjälte ! 
Du är Neapels nya Munaciello ! 
Kan du simma ? 
Jag ligger på nivå åtta . 
Åtta ? Snart blir det nivå nio . 
Vart är du på väg i de där kläderna ? 
- Jag ska ta en promenad . 
- Så här sent ? 
- Vad ska du med skateboarden till ? - Inget ! 
Vad har du där för något ? 
Stal du och dina vänner statyetten ? 
- Sasà ! 
Enzo ? 
- Trodde du att du kunde lura mig ? 
- Jag ? 
Vad menar du ? 
Du var den enda som kände till statyetten . 
Du bad killen på skateboard att stjäla den och lagfarten , eller hur ? 
Vad pratar du om , Enzo ? 
Slyngeln slängde sig ner i brunnen utanför Palazzo Spinelli . Han föll pladask och statyetten med . 
Er plan har gått i stöpet . 
Skulle jag ha en plan ? 
Ser du inte att jag inte är en enda röra ? 
Vet du vad ? 
Imorgon ska du hämta statyetten . 
Annars kommer jag se till att du får det ännu värre ställt . 
Är det uppfattat ? 
Javisst , Enzo . 
Vad vill ni ? 
Vår vän dök ner i havet och vi hittar honom inte . 
Du måste hjälpa oss ! 
Vi vet att han lever . 
Han tog sig in under marken för att hitta Wonderboy . Han stal en statyett från vår hyresvärd . 
Vem letar han efter ? 
Wonderboy . 
Han är ungefär som Munaciello . 
Varför skulle han bry sig om Munaciello ? 
- Jag förklarade bara . 
- Munaciello har alltid funnits . 
Det är folket ... som har glömt av att staden är full av magi . 
Men nu måste vi möta honom . 
Hur tar man sig ner dit ? 
Det kommer inte att bli enkelt . 
Kom här . 
Den enda vägen in ... går genom Gaiola . 
Det är den mest hemsökta platsen i hela Neapel . 
Naturligtvis . Vi måste till den hemsökta ön . 
Rafè , vi måste hitta vår vän . Håll tyst nu . 
Jag vill hellre prata , annars blir jag nervös . 
Titta ... Vem vet hur många spöken som finns där . 
Vad är det där ? Båten rör på sig av sig själv ! 
Hörni , det är jag som drar hit den . 
- Hoppa på . 
- Han är helt från vettet . 
Kom igen . 
Sasà ! 
Är det du ? 
Sasà är inte tillbaka än . Han lämnade sin mobil på sitt rum . 
Han är säkert med sina vänner . 
Antò , vart ska du ? 
Vad pågår egentligen ? 
Francè , ursäkta . Är Gennaro och Raffaele hemma ? 
Ja , de sover . 
Vi åker till Brescia imorgon . 
- Vart ska hyresvärden ? 
- Antò , vad ville du ? 
Oscar ! 
Antò , kan du berätta vad som händer ? 
Jag måste låna din scooter . Jag ska följa efter hyresvärden . 
Vill ni verkligen gå ner där ? 
Det är okänt område . 
Vi tar livet av honom . 
- Bra tänkt . Det gör vi . - Nej ! Vänta ! 
Det lär finnas en annan väg in . 
Men ingen har faktiskt använt den . 
Nu artar han sig . 
- Vissa delar har rasat in . 
- Var är det ? 
På Gaiola . 
Du är galen . 
Det spökar på Gaiola . 
Ja , därför ni borde ge upp . 
Gennà , det finns ingen mottagning här . 
Vi är under marknivå , vad trodde du ? 
Jag tror att jag ser en stege . 
Det är precis som Clemente sa . 
Ja . Vi får hoppas att han hade fel om resten han sa . 
Fortsätt . 
Gennà ! 
Jag hatar det här stället . 
Vad hände ? 
Det var inget , Rafè . Det var bara vinden . 
Det här är Sasàs . 
Vi måste skynda oss . 
Alfrè ! 
Angelica ! 
Ja Angè ! 
Inne i statyetten finns det en skattkarta . 
Det var längesen vi sågs . 
Letar du efter statyetten ännu ? 
Har du inte fått nog efter allt som har hänt ? 
Hur kan jag ha fått nog om det inte är över än ? 
Vet du vad hyresvärden letar efter ? 
Det är en statyett , men jag vet inte varför . 
Jag är säker på att ungarna är involverade . 
En gorgon ... 
Terè ? 
Vilket ställe ... Nu går vi härifrån ! 
Vi måste hitta honom . 
Var inte dum , Rafè . 
Vi ska träffa Clemente om två timmar . 
Vad är du rädd för ? 
Ingången måste vara här . 
Terè , vart ska du ? 
- Vad gör du ? - Terè . 
Terè ... 
Vad gör du ? 
Teresa ! - Teresa ! - Teresa ! 
Kom igen . 
- Tonì ? 
- Vad ? 
Går vi verkligen uppåt ? 
Hur vet du vilken väg vi tar ? 
Prata mindre och knata mer . 
Annars funkar inte mina superkrafter . 
- Hörde du det ? 
- Ja . 
Det här är avloppet . Jag tror att vi närmar oss . Följ mig . 
Kom . Var inte orolig . 
Teresa ! 
Jag ser inte ett dugg . 
Kom hit , hörni ! 
Vad gör vi nu ? 
Vad tror du ? Vi går efter . 
Sasà , släng ner den . 
Vi kommer , Wonderboy ! 
- Terè ! - Teresa ! Teresa ! 
Kom här , hörni ! 
Kom hit . 
- Aniè ! 
- Hörni ! 
- Aniello ! - Aniello ! 
Aniè , vi hittade dig ! 
Kom här . 
Jag visste att ni aldrig skulle lämna mig ! 
Hörni , vi var inte galna . 
Wonderboy finns på riktigt . 
Titta ! Han är Munaciellos efterträdare . 
Han stal statyetten från hyresvärdinnan ! 
Vi gjorde det ! 
- Hurra ! - Jag har saknat er ! 
Vi saknade dig med . 
Han är borta ! 
Och nu då ? 
