Hej , Crayola . Gul ? 
Gul som solen , gul som en anka . 
Utmärkt val . Alla älskar ankor . 
Okej , gör orange . 
Vit . 
Grå . 
Svart . 
Beige . 
Tack . Men jag är här för att jag var vaken hela natten och tänkte på att ni måste tillverka en genomskinlig krita . - Genomskinlig ? - Ja , som färgen . 
Men genomskinlig är inte en färg . 
Vad kallar du det här då ? 
- Vad då ? 
- Det känslomässiga utrymmet . 
- Men ... om kritan är av genomskinligt vax och den inte lämnar synlig färg , - vad är poängen ? - Det är omöjligt ! Varför gör du det här ? 
- Varför behöver du den ? 
- Den finns redan . 
Se på vattenglaset . Det är helt klart genomskinligt . 
Vissa saker är inte normalfärg eller följer regnbågens regler . 
Tänk på luft , dofter eller minnen . 
Borde inte de få ha egna färger ? 
Att färga nåt genomskinligt visar att saker och ting är olika och det är okej . 
Att färga nåt genomskinligt förändrar våra föreställningar om färgläggning . 
Tack för att du kom förbi . Du har gett oss mycket att tänka på . 
Om vi går vidare med genomskinliga kritan , vad ska vi kalla den ? 
Kalla det fantasmas . 
- Fantasmas ? - Det betyder spöken . 
Varför plural ? Varför inte fantasma ? 
Det heter blå , inte blåa . 
För att jag gillar det . 
Javisst . Men logiskt sett borde det vara fantasma . 
Du har nog rätt . 
Kalla det fantasma . Singular . Inget " s " . - Bra . - Bra . 
Var är min bil ? Där är min skjuts ! 
Hej , är du Julio ? 
Välkommen till Chesters . 
Bara några grejer . 
Stäng dörren försiktigt , avinstallera din Uber-app och ladda ner Chester . Det är den enda app som du kommer att använda . 
CHESTERS BIL Vad är en Chester-app ? 
Chester är helt enkelt ett alternativ till Uber men alla intäkter går till Chester . 
Du kan boka skjuts med mig via appen och få tillgång till forumet där användare delar med sig toakoder för olika Chipotle-restauranger . 
Vi jobbar på gräsrotsnivå . 
Och om du är en äldre medlem så kan du bli upplockad och avsläppt även om jag redan har en kund . 
Teven måste vara på hela tiden och endast spela Melf . 
En till dig och en till dig . 
Hur bär du dig åt ? 
Grace , akta dig . 
Vad är du för nåt ? 
Jag heter Melf och kommer från planeten Melf . 
Snälla , kan vi behålla honom ? 
Okej . 
Melf älskar kakor och spagetti . 
Jeff ? 
Jag hörde ljud på nedervåningen och trodde att det var tjuvar . Det visade sig bara vara Melf som äter kvällsmål alldeles ensam . 
Hjälp mig att städa undan det här . Inga ursäkter , Melf . 
Vet du vad ? Lägg dig igen . - Jag kan städa undan . - Okej . Godnatt . Stanna inte uppe för länge . 
Vi måste vara försiktiga , Melf . 
Mel älskar kakor ... och spagetti . Och Jeff . 
Jeff gillar Melf med . 
Melf vill inte vara utanför . Melf vill vara först . 
När ska Jeff berätta för Nancy om Melf ? 
Snart . 
Jag älskar dig . 
Ni skrämde mig ! Vad håller ni ... ? Vad håller ni ... ? Lyssna ... 
Vad fan pratar du om ? 
- Skämtar du med mig ? - Okej . Ut ! Stick , Jeff ! 
SJUTTON ÅR SENARE ... - Hej , pappa . - Hej , älskling . - Hej . 
- Hej . - Får jag komma in ? - Självklart . 
Tack för inbjudan . 
Jag blev förvånad att du ringde , Grace . Jag heter Toast nu . Ja . 
Din mamma dog och gav dig ringen . 
Jag skojar . Åh , herregud . Min lilla ... - Toast . - Toast ska gifta sig . 
- Du kommer att gilla henne . 
- Henne ? 
Skojar du ? Förlåt , jag ... Din styv-Melf kommer att bli så glad . - Pappa . - Har ni en bröllopsönskelista ? 
- Vad du än vill ha så köper vi det . - Jag vill inte ha Melf på bröllopet . 
Jeff , du kan inte gissa vem jag stötte på i affären idag . Jag ... 
Jeff , Melf lämnade några varor i bilen . 
- Jag kan hämta dem . - Vänta , pappa . - Pappa . - Är du hungrig ? 
Jag skulle precis gå . 
- Låt Melf fixa lite mat . 
- Jag måste verkligen gå . 
Hur vore det med lite kakor och spagetti ? 
Julio ? - Julio ? 
- Där är Bibo . 
Lägg av . Är det din assistent ? Ja , som en sekreterare . 
Hej , Bibo . 
- Välkommen till Chesters , Bibo . 
- Tack . 
Jag behöver ta ledigt imorgon för att rengöra tänderna . 
- Men du har inga tänder . 
- Det står i kalendern . 
Ja , men du har inga tänder . 
Jag har en kupong . Jag vet . Lyssna , det är helt okej att du tar ledigt imorgon . Det är helt okej att du går till tandläkaren . Men jag vill inte att du går dit och blir besviken när det inte finns nåt att bleka . Manipulatör . Jag vill ha löneförhöjning . 
Har du några ärenden som inte har att göra med Bibo ? 
I själva verket så fick du ett sånt här . BRÅDSKANDE 
Det verkar vara brådskande . 
Julio , du ignorerar det igen . Breven bara växer på hög . 
De är troligen från din hyresvärd . 
Vad är det för lockrop ? 
Julio , dagdröm inte . 
Hör ni det ? - Hör ni det ? - Nej . Vad då ? 
- Jag hoppar ut här . - Okej . 
- Trevligt att träffas , Chester . - Detsamma . Ha en fin dag . 
Du med . 
Hej . Vad är det här ? 
Vad är det för ljud ? 
Det är ett litet ostron med små diamanter . 
Det är unikt . Sällsynt . Vackert . 
Jag tar det . 
- Vad då ? - Leverfläcken bakom ditt öra . 
Den ser ut som ostronets skugga . 
Det är inte en leverfläck . Det är ett födelsemärke . 
Jag har kollat upp det . 
Det är precis samma storlek . Så ... 
Så konstigt . 
Hon sa att det var en förbannad antikvitet , så jag måste köpa den . Perfekt . Den är perfekt . Den ende i sitt slag . Tack . 
Åh , herregud . Som hans lägenhet . Har du sett den ? 
Den är jättefin . 
Det här kommer att bli en stor grej för dig . 
Jag tappade den . 
- Nej . - Ja . 
- Ostronet ? 
- Ja . Nej . 
- Hittade du det ? 
- Nej . 
Jag vill sticka . Vill du dela en Chester med mig ? - En vad då ? 
- Chester . 
Okej . Är ni redo ? Jag ska först släppa av Amina eftersom hon är lärare , men ni står näst på tur . 
Åh ! Där är byggnaden som jag ansöker till . 
Ska du flytta in i Capital Ones bostäder ? 
Exxon Mobils bostäder . 
Julio , de har en simbassäng . 
Jag har hört att det är fint . 
- Men visst ber de om den där grejen ? 
- Bevis på existens ? 
Ja . De ber om det för alla lägenheter nu . 
Jag bryr mig inte om nåt jäkla bevis på existens . 
Jag behöver inget bevis . 
Uber försökte skaffa ett åt mig . Jag sa : " Ni vill ta hälften av de pengar som jag tjänar och ta betalt för ett ID som bevisar att jag existerar ? " Jag existerar . 
Bra . 
Jag har inget bevis och vill inte ha det . - Jag vill inte ha det . - Såja . Släpp ut det . 
Jag ser hemsk ut på mitt bevis . 
EXISTENSBEVIS - Vad jobbar du med , Vanesja ? 
- Det uttalas Vanessa . 
J:et är tyst , som en giftig blomma . 
Oj . Jag är en mycket viktig talangscout på ett mycket viktigt uppdrag . 
Hon är en skådespelare som låtsas vara min agent , men hon har gjort det så länge att hon nu gör vanliga scout-grejer . 
Det är lite oklart . 
Vänta lite , anlitade du en agent för ditt bevis ? 
- Inga fler frågor , Chester . 
- Så hemlighetsfull . 
Du då , Julio ? Vad sysslar du med ? 
Julio träffades av blixten som barn . 
Ända sen dess har hans syn på världen varit lite annorlunda . 
När jag vaknade fick jag ett intyg på att skippa gym för resten av livet . 
BARNLÄKARE Jag laminerade det och visar det när folk ber om bevis . Okej . Förresten , vad gjorde du i skogen ? 
Jag minns inte . - Han bajsade . 
- Det spelar nog ingen roll . 
Han torkade sig när blixten träffade . 
Men han utelämnar det från historien på grund av skamkänslor . 
Men vad gör du ? 
Jag är lärare . - Du är ... - En Julio . 
Det är vad han gör . 
Förklara . 
Jag vaknar och bara är en Julio . 
Det är fantastiskt . Idag konsulterade han för Crayola och imorgon har han ett möte med NASA för att döpa om en konstellation . 
Jag kan känna det inre livet hos former , färger , ljud , nummer och bokstäver . Jag började nyss med bokstäver . 
Låt mig ge er ett exempel . 
Ni vet hur bokstaven Q är placerad alldeles för tidigt i alfabetet ? 
Vad menar du ? 
Den borde vara med de andra avantgardebokstäverna . X , Y och Z. Q bad inte om att vara tidigare . Föreställ er hur det skulle kännas . 
Förtjusande . Så trevligt och lätt . Ge en applåd för P. 
Och nu en applåd för Q. 
Alla bokstäver har varit så tillgängliga tills Q intar scenen . 
Hej , jag är Q. 
Ni kommer alla att dö ! Jag vet inte varför ! Era jävlar . 
Tack . 
Nästa sång heter : " Din gylf är öppen och din kuk hänger ut . " 
Ingen förstår honom . Q är för tidig i alfabetet . Lägg av , jag sitter i kläm mellan dessa två ... normisar . 
Förlåt , men det är vad de är . 
Vem fan har du på scenen nu ? R. 
Lyssna på honom . De slukar honom . 
Jag är inte lika lättbegriplig . 
Därför måste du lägga mig sent . När alla är fulla . - Vi har pratat om det . 
- Jag bestämmer inte ordningen . Vet du vad ? 
Den här klubben suger och du med . Jag är stolt över min nisch . Jag bryr mig inte . 
Jag skojar bara . Kom igen . Du känner mig . Ge mig en chans . 
Men Q fortsätter att vara Q. 
Social trygghet Åh , du förfaller Din pensionsplan är inte okej Ha en bra dag - Så fantastiskt . Vad är det ? - Hörru ! Kom igen . 
Trevligt att träffas . Jag är O. Vet du vad som är skillnaden mellan dig och mig ? Vad då ? 
Din pinne . 
Ta bort den . 
- Ja , men då skulle jag vara ... - Jag . 
Min inhoppare . 
Jag har så många spelningar . Orange , orangutang , ollon . Jag är två gånger i det ordet . 
Lyssna , jag har fullt upp . Jag behöver extra hjälp . Ring mig när du inte längre vill vara en arbetslös bokstav . 
Jag kan också göra så . 
Ingen köper det Q säljer . Det finns ingen marknad för udda . 
I flera år måste Q hitta på andra sätt att betala räkningarna . POPNYHETER Medan alla konventionella bokstäver badade i möjligheter . 
... blir den populäraste konsonanten i alfabetet . 
F gör sig redo att skriva under ett kontrakt värt flera miljoner för att börja ett nytt ord med Amerikas älskling , bokstaven B. 
Sen hände det värsta . Udda blev plötsligt coolt . 
Vi är W , X , Y och Z. Vi följer inte dumma regler och vi är inte snälla . 
Och Q missade tåget . 
Ni har aldrig sett nåt liknande . Vi krossar reglerna , vi ställer oss inte i kö ... 
Orättvisan blev allt mer uppenbar vilket snart blev för mycket för Q. 
Under alla år som han ägnade sig åt sin konst . CBGB PRESENTERAR " Q " MED V CBGB PRESENTERAR Q MED W OCH SV Han känner sig fången och bestämmer sig för att bryta sig loss . 
Fan ! 
Okej , så hyser nån av de konventionella bokstäverna i alfabetet agg mot er ? 
Tja , bokstaven G har skickat meddelanden till oss . 
- Hallå ? - Hej . - Hej , det är Q. 
- Jag vill bara säga en sak . Vi skulle nog inte vara här utan Q:s inflytande . 
Jag känner dig inte men ... Hans verk har påverkat mig och jag talar nog för oss alla att vi inte hade varit här om inte Q hade tänjt på gränserna . Han var inte ute efter berömmelse eller ära utan det obevekliga , orubbliga engagemanget för äkthet . Q gjorde publiken obekväm långt innan udda var coolt . 
Ser du detta så ska du veta att jag är ett stort fan . 
Är du där ? Hallå ? Dra åt helvete . 
Visst kände ni det ? 
Allt detta bara från att se på bokstaven Q ? - Jag sa ju , det är vad jag gör . 
- Ring mig om du vill boka honom . Så fixar Vanesja det direkt . Amina , vi är framme . Amina . 
Förlåt . Tack . Hejdå . 
Jag kan inte sluta tänka på den . 
Jag såg den för en vecka sen . 
Det var sent och jag var en av de få kvar i skolan . 
DAMERNAS UR BRUK Medan jag hängde över toalettstolen funderade jag på teckningarna som pojkarna hade gjort i båset . 
Sen ... såg jag den . I hörnet av båset , som om den gömde sig från sina vänner , fanns en penis med sitt huvud bortvänt från betraktaren . 
Vad kan den betyda ? 
Var kuken ledsen ? 
Är den förkrossad över alla förväntningar om manlighet ? 
Eller levde den bara sitt eget liv ? 
Jag kunde inte ignorera detta . 
Jag måste veta vem som tecknat den . 
Det kanske var en av bögarna ? Nej . Bögar tecknar inte penisar . De tecknar ögon . 
Med långa , läckra ögonfransar . 
Vänta lite . 
Läget , Rick ? 
På pojkarnas toa , tecknade du en penis som undviker betraktarens blick ? Så här ? 
Varför har du på dig en lila tröja ? 
Lila är en tjejfärg . Du ska inte ha på dig det . 
Lägg av . 
Han ska inte ha på sig det . 
- Varför inte ? 
- Din subba . 
Okej , kvarsittning . 
Jäkla mobbare . 
Michael ? 
Har du ritat den här ? Ja , för att jag är kille , din subba . 
Michael . Varför ser penisen ut så ? 
Ibland så ... känns det att som kille finns det saker jag inte kan göra . 
När jag ser killar göra saker som att ha på sig lila kläder så blir jag arg . 
Så jag sparkar dem för att påminna dem om reglerna . 
Du ser mig vara taskig men ... jag är taskig för att du ska se mig . 
I själva verket ... så ser ingen mig . 
Fröken Roberts ... jag är fången . 
Jäklar , fröken Robert . Du är gift ! 
Subban är så jäkla kåt . Jag svär . 
Vad är det här ? 
- Var går de här nycklarna ? 
Jag och grabbarna var fulla igår och hittade dem vid ett staket . 
Vad ? 
De var nog där så att nån skulle hitta dem . 
- För att ta sig in nånstans ? - Ja . Nu är de utelåsta . 
I brevet står det : " Gracias , mama . " 
Nu blev nån dam som du inte känner utelåst sent igår kväll . 
Är du arg på mig ? Nej , jag är inte arg . Jag är bara ... Jag är bara förbryllad . Till och med min flickvän hatar mig . 
Jag blev inte befordrad . Hallå ? Jag behövde lätta på trycket med grabbarna . 
Jag måste be dem att komma ut eftersom jag inte är Jared . 
När Jared skickar meddelande till gruppen så är alla redo . 
Det är dödstyst när jag gör det . 
När jag äntligen har lite kul och gör ett litet spratt så får du mig att må dåligt . 
Vill du se True Women of New York ? 
Är du säker ? 
Vänta . 
Ja , men du måste ge den tillbaka , för den måste ges till forskarna . DRÖMANALYS-KIT 
Det sägs att svaren till alla våra problem finns gömda i våra drömmar . 
Julio , rullar du fortfarande ? 
Nej , det gör jag inte . Det där var högst opassande . 
Hämta din gummianka . Dags för vår dusch . 
Vår vadå ? 
Ibland känns det som att jag inte känner dig . 
Hej , hallå . 
Jag har haft en återkommande dröm . 
Jag är i ett rum . Jag har på mig en hög strutmössa . 
Plagget är gjort av silke eller bomullsblandning , det kvittar . 
Jag sitter vid en nån slags manick . Väldigt genialisk , faktiskt . Den låter mig läsa utan att behöva vända sida . Fattar du hur irriterande det är att spela in en dröm 
- medan du lyssnar på det där ? - Skrik inte på mig . 
Förlåt , det var inte meningen att skrika . Det är lugnt . 
Manicken låter mig läsa en hel bok utan att behöva vända sida . Men sen känns det lite varmt så jag vill öppna ett fönster . 
Men jag går till fönstret och det leder ingenstans . 
Jag öppnar nästa fönster . 
Samma sak . 
Och igen . Jag går till nästa fönster och samma sak . 
Jag öppnar dörren och inte heller den leder nånstans . 
Sen ser jag en dörr tvärs över rummet . 
Den leder ut . Det snöar . 
Folk går omkring i uniform i såna här alldagliga svarta pufferjackor . 
Om jag går ut måste jag ta på mig en för att hålla mig varm . 
Sen ser jag den . En svart pufferjacka med mitt namn som kallar på mig och säger : 
Jag återvänder till rummet , skräckslagen . Rummet håller på att krympa , så jag försöker lämna rummet men jag kan inte på grund av min stora , vackra hatt . 
Enda sättet att lämna rummet är genom att kompromissa , men hur ? Sen vaknar jag och drömmen är slut . 
- Ett till har anlänt . - Ett till vad då ? 
Lägg det med resten . 
Det ser inte viktigt ut . 
Det är från din ... hyresvärd . 
- Läser du min post ? - Med min röntgensyn . Jag öppnade inte det så det är inte ett brott . Det är mycket viktigt . 
Ser det här födelsemärket större ut ? Jag tycker det . 
Jag oroade mig inte över det men Chester sa : " Det ser illa ut . Du borde kolla upp det . " 
Borde jag kolla upp det ? Om du är orolig så borde du kolla upp det . 
Du skulle ha sett deras ansikten . De sa : " Herregud , " och deras hakor föll ner till golvet . 
Det står att du måste flytta . 
De gör om byggnaden till ett General Mills-kafé och bostäder . 
Jag borde gå till läkaren . 
Julio , du behöver en ny lägenhet . För att få en ny lägenhet behöver du bevis på existens . 
Nej , jag kan inte tänka på lägenheten eftersom jag är sjuk . 
Nej , Julio . Försvinn inte i dina tankar . 
Kom tillbaka . Bemöt det verkliga problemet . 
Den har nog växt . Den har växt . Den har definitivt växt . 
Åh , herregud , det här blir jobbigt . 
