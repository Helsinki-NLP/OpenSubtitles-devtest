Vi har listat ut det ! I TIDIGARE AVSNITT Fotot är en ledtråd ! 
En mor gör allt för sina barn ! 
Jag är ingen mor ! 
Om Clemente hoppade ända däruppifrån , så har havet ha tagit honom . 
Oroa dig inte , donna Angè . 
- Jag fixar det här . 
- Nej ! 
Hörde du inte vad hon sa ? 
Du är inte boss längre . 
Fotot inuti statyetten togs på Arkeologiska museet . 
Om jag kan väcka elixiret till liv , kan jag kanske träffa mamma igen . 
Antò ? Hör du mig ? 
Hans gömställe ... 
Hon ville gå till katakomberna med prinsens elixir . 
Den farligaste delen är precis ... 
Det här är alla Munaciellis gömställe . 
Vi önskar er en trevlig kväll . Utgången är här borta . 
Utgången är härborta . Tack så mycket . 
Vi önskar er en trevlig kväll . 
Tack så mycket . 
- Adjö och tack . - Ursäkta ! 
Utgången är hitåt . 
Nu stänger vi . Tack för ert besök . Hej då . Adjö . Ha det så fint ! 
Nu är det dags för middag . 
- Vad är det där ? Hördu , Savè ? - Vad ? 
Ser du ljuset och röken därborta ? 
Vad är det för nåt ? Spökglober ? 
- Vad ? 
- Spökglober ? 
- Ja , säkert . Det heter " ljusklot " ! 
Ta en kaffe från automaten . 
Men gör det fort . Jag ska låsa porten . Oroa dig inte . 
Det är en underlig känsla ikväll . 
Sankt Sasà åstadkommer mirakel ! 
Det är inget mirakel . Det här är en cykelgenerator . 
Titta här , Rafè ! 
Här står namnen på alla Munacielli . 
Sabello . 
Lucio . 
Silvestro . 
Alfredo ! 
Han är den sista ! 
Det här är på riktigt , hörni . 
Vi är i Munacielli-gömstället . 
Det måste ha varit Alfredos ande . Han ledde oss hit med hjälp av Genuasås . 
Det var här han gjorde Maradonastatyetten . 
Det här måste ha varit hans verkstad . 
- Titta där ! 
- Vad är det ? 
Vem hade väntat sig det här ? 
Han sparade alla artiklar om honom . 
" En figur från en julkrubba hittades inuti ett vitrinskåp där en värdefull klocka tidigare hade haft sin plats . 
Vår stad anser honom inte vara nån tjuv , utan en modern Robin Hood , som stjäl från de rika och ger åt de fattiga . " 
Du ... Hur mår du ? 
Jag känner mig bättre . 
Teresa har varit här . 
Vi måste hitta henne . 
Först måste vi hitta Clemente . 
Försiktigt . 
Donna Angè , vad händer ? 
Det var 25 år sen sist . 
God kväll . 
Vi stänger nu , tyvärr . 
Det är akut . Vi måste komma in . 
" Akut " ? Hur menar ni ? 
Det går inte ikväll . Snart kommer våra tekniker De ska installera en ny utställning : " Parthenope - Neapels sång . " 
Jag lämnar en donation . 
En donation . 
Var god , stig på . 
- Ta hand om det . 
- Vänta . Donationen . 
Tusan också . 
Den här vägen , tack . 
Välkomna . 
Ni är tre stycken . 
Jag kan tända för er . 
De måste ha gått in genom den andra ingången . 
Jag skulle absolut ha märkt om en grupp barn var kvar på museet . 
Vad gör vi nu ? 
Här . Varsågod . 
Barnen har länkat sina mobiler till datorn . 
Nu ska vi bara spåra dem , så ser vi var de är nånstans . 
- Lösenordet ... 
Jag kanske stavade fel . 
Lösenordet har alltid varit " Kom igen , Neapel . " 
- Vi valde det alla tre ihop . 
- Jag visste det . 
De är inga småglin längre , Mariù . 
" Ingen ser honom som tjuv . 
Han är bara den senaste Munaciello . " 
Det var en fin historia om Munaciello , men vad gör vi nu ? 
Titta här , hörni ! Kom ! 
Vad är det här för ställe ? 
Det är ett mörkrum där man kan framkalla foton . 
Det här är negativet för samma foto som fanns inuti statyetten . 
Får jag se . 
- Otroligt ! 
- Det måste vara en annan skattkarta ! 
Men hur framkallar man fotografier ? 
Vi behöver en tutorial-video . 
Har du nåt nätverk här ? 
Mobilen fungerar inte härnere . 
Etthundratjugosju aviseringar ! 
- Oj , de måste vara jätteoroliga . 
- Än sen ? 
Vi måste hitta skatten . Annars var allt det här förgäves . 
Nej , vi måste hitta Teresa ! 
Har du glömt det ? 
Hon skulle inte ha stuckit ! Sluta bråka ! 
Hörni , om vi lägger ner nu , så skulle allt vi gjort vara förgäves . 
Vi framkallar fotona . Vi ringer upp föräldrarna och letar efter Teresa . 
Ge mig din telefon . Vi måste hitta en tutorial . 
- Salen är därborta . 
- Det var på tiden ! 
Jag är redan stressad av att hinna med allt på en kväll . 
Vi behöver inga förseningar . 
God afton . 
Var försiktig ! Sirenens dräkt är jättedyr ! 
De har till och med lämnat fotavtryck . Hur har ni inte sett det ? 
Vad är ni för vakter ? 
Clemè . 
Nu får du göra din del av avtalet . 
Spåra dem . 
Tonino ? 
Det är jag , Clemente ! 
Kom igen ! 
Det här är ingen lek . 
Du kan lita på mig . 
Jag hade rätt . Ni känner varandra . 
Sänk rösten , annars hittar de oss . 
- Du ljög . 
- Antò . 
Där är han ! 
Vad händer nu ? 
- Antò . De kommer att hitta oss . - Släpp mig . 
Ande , vars hjälp jag ber om . Jag har en gåva till dig . 
Det är ingen juvel . Det är något ännu mer värdefullt . 
Det är ett elixir som för döda tillbaka till livet . 
Jag trodde att det var det här du ville . 
A mortis limine restituo . 
Mamma ? 
Såg du ? Jag gav elixiret till anden så att du kunde komma tillbaka . 
Du var jätteduktig . Men jag har aldrig lämnat dig . 
De döda lämnar en aldrig . 
Alla fina saker som vi varit med om , alla fina minnen och de dåliga ... De blir en del av dig . 
Döden kan aldrig utplåna dem . 
Jag vill ha dig hos mig igen . Jag vill att du gör min skollunch . Jag vill att du ska borsta mitt hår varje morgon . 
Du lät mig aldrig borsta håret , Terè . 
Vill du veta vad hemligheten var som gömdes i ampullen ? 
Du skulle fylla den med tre ting . 
Rädsla , kärlek och smärta . 
Dessa tre ting är vad livet handlar om . 
Nu har du lärt dig det här och kan återgå till att leva utan att vara rädd att få lida . Och även om jag inte är kvar , så har du dina vänner , din morbror och din pojkvän . 
Men jag kan inte leva utan dig . 
Farväl , mamma . 
Jag älskar dig . 
Kul att han känner sina barn så väl . 
Vi har hållit på med det här i tre timmar . 
Jag känner mina barn , ska du få se . 
Jag har listat ut lösenordet . 
" Jag hatar Brescia . " Jag lägger till ett utropstecken också . 
Bra jobbat . 
Nu när du har visat att du inte känner dem kan jag gå till polisen . 
Terè ? 
- Antò ? - Låt mig vara , Tonì . 
Snälla , lyssna på mig . 
Om det blir känt att vi känner varann , kommer du också att råka illa ut . 
Det är bäst så här . 
Lita på mig . 
Okej . 
Men få mig inte att se ut som en idiot . 
Tonì , titta där . 
Vi hittade dem . 
De liknar grenar . Men de är tunnlar . Ge mig fotot . 
Nu får du lita på mig . 
Du är ett geni , Antò . 
Men hur ska vi kopiera det ? 
- Kan vi använda den där ? 
- Vänta . 
Jag går . 
Äntligen hittade jag dig . 
Ursäkta mig ? 
- Vad vill du ? - Varsågod . Här får du till kaffe . 
Stick härifrån ! 
" Här får du till kaffe . " 
Fy , vad det stinker ! 
Ingenting stoppar Capuozzo Enzo ! 
Gennà , titta på den här antikviteten ! 
Den är trasig . 
Det kokar ! 
Jag är så hungrig . 
Jag vill lägga en liten tomat där . 
Ska vi inte koka lite pasta sen ? 
Vilka är ni ? 
Är ni de där försvunna odågorna ? 
Var är statyetten ? 
- Och vem är du ? 
- Jag är gubben som ska klå upp er . 
Statyetten . 
Vad var det inuti ? 
Nu har jag fått nog , okej ? 
Du har rätt . 
Det låg en skattkista inuti statyetten , men Tonino tog den ! 
- Och nu är vi fast härnere ! 
- Vet du vad vi ska göra ? 
Nu ska vi alla , lugnt och fint , leta upp Tonino . 
Annars kommer det att bli obehagligt ! Jätteobehagligt ! 
Vad skulle ni göra , ta en tur i underjorden ? 
- Vi måste få ut dem därifrån . 
- Ja . 
Men vi har fastnat här . Titta . 
Sista frågan vi ska besvara är deras favoritlåt . 
Vilken då ? 
Säkerhetsfrågorna ... 
Vi kan inte lösenordet . 
- " Gaiola ger oss lycka . " - Nej ... 
- Okej ! 
- Bra jobbat , Teresa ! 
Utmärkt . 
- Det står att de är här . 
- Men var ? 
Kanske är det där ? 
Vänta på mig här . 
Det är trångt , men jag slinker igenom . 
Var försiktig . Det är farligt . 
Hon vet vad hon gör . 
Var försiktig , Terè ! 
Den här stan är magisk . 
Du knockade mig nästan när vi först träffades . 
Och nu tänker jag kyssa dig . 
Tonì . 
Din tid är nästan ut . 
Ge upp . 
Därborta ! 
Det är radion som de stal från mig . 
- Vi delar på oss . 
- För dem till mig ! 
Ge mig ett stort leende . 
Du är så vacker . 
Vad är det , Angè ? 
Alfredo . 
Alfredo ? 
Vad har han med den att göra ? 
Det är som att han försöker säga nåt till mig . 
Jag går ! Vänta ! Jag hörde nåt . 
Titta , Antò . 
" Zeus var så svartsjuk att han höll på att tappa vettet . 
Han kunde inte acceptera att sirenen Parthenope var förälskad i kentauren Vesuvius . " 
Se in i varandras ögon , seså ! 
Bra . 
De här två blir perfekt . 
Ring dansarna . 
Ge dem en ursäkt . Säg att tillställningen är uppskjuten . Seså . 
Spela musiken som jag bad om . 
Vad är det för musik ? 
Vilka är ni ? 
- Ursäkta oss ett ögonblick . 
- Vad menar ni ? 
- Vi arbetar ! 
- Ta det lugnt ! 
Din läspande byracka . 
Ni är de sista vi behöver ! 
Såg de att det är vi ? 
Nej , men hyresvärdinnan är distraherad . 
Det här är vår chans att fly . 
Sätt fart . Jag vill se om det är farligt . 
Jag måste gå samma väg i så fall . Kom igen ! 
- Det här är giftig gas ! 
- Sätt fart ! 
Jag sparkar skiten ur er ! 
Sätt fart ! Nu kommer jag ! 
Vad gör ni ? 
Låt mig se . 
Vad är det där ? 
Det är sirenen Parthenope . 
Om man hör hennes röst , så dör man strax . 
Nej . 
Jag kan inte dö . Inte nu . 
Nej . 
- Spring , hörni ! 
- Vänta på mig ! 
Den här vägen , hörni ! 
Jag visste att det var du ! 
Terè . 
Ingen kan stoppa oss ! 
Kom nu . 
Hur är det med dig , Clemè ? 
- Jag är okej . 
- Vad hände ? 
Ingenting . Det är okej . 
Nå ? 
- Vad är det här ? 
- Ingenting . 
Du behåller den här . 
Innan vi går till underjorden måste jag hämta nåt jag behöver . 
Vi ses vid min husbil . 
- Berätta vad som pågår . 
- Det är inget , Antò . 
Jag möter Clemente , sen går vi och hittar skatten och barnen . 
- Men det är för farligt ... - " För en kvinna " ? 
Jag räddade faktiskt livet på dig ! 
Clemente ? Var är Clemente ? 
Han har rymt igen ! 
Stick efter honom ! 
Sluta ! 
Donna Angè , vi har gjort allt vi kunde ! 
Om du inte har pengar får du inga mannar . 
Hur vågar du ... 
Jag fick betala donationen för att komma in ! 
Chihuahua gjorde rätt som lämnade dig . 
Kom . Vi drar . 
Tölpar ! 
Ni ska få betala för det här ! 
Era fähundar ... 
Varsågod . 
Den här låg i statyetten . 
Du förstörde våra liv för ett litet foto . 
Angè , jag har gömt skattkartan i den här statyetten . 
- Om nåt skulle hända mig ... - Varför skulle nåt hända dig ? 
Om något allvarlig händer , måste du komma och hämta mig . 
Jag är höggravid ! 
Gå inte . 
Skit i skatten . Jag vill ha dig . 
Jag vill att vårt barn ska ha en far . 
En far som dina föräldrar inte accepterar ! 
Jag vill inte vara osynlig ! 
- Vi sticker ! 
- Vart ? 
Jag vet inte vart ! 
Men vi rymmer tillsammans ! 
- Du fattar inte . 
- Vad är det jag inte fattar ? 
Folk här ser på mig som en tjuv . 
Jag är trött på det . 
När jag hittar Lautrecs skatt , blir jag Neapels nya hjälte . 
Fattar du , Angè ? 
Neapels nya hjälte , älskling . 
Jag hoppas att du blir det . 
Jag vill inte delta i din galenskap . 
Kan du stanna här hemma en stund ? 
- Ja . 
- Jag ska leta efter din syster . 
Jag trodde aldrig att du skulle rädda mig . 
Du bäst , pappa . 
Trodde du att jag bara skulle ge upp ? 
Ja . 
Du är väl okej ? 
Nu är allt bra . 
Det är bra . Precis som vanligt ... 
Jag gör alltid grejer för andra . Varför ? 
Vad hände med Tonino ? 
Han gick till Clementes husbil . De ska leta efter skatten . 
Han brydde sig aldrig om oss . 
