Alice , älskling , prata med mig . 
Du måste hålla dig vaken . Du får inte somna . Alice ! 
Hur hamnade du där ? 
Alice ? Älskling ? Min älskling . 
Är du ett spöke ? 
Mamma är strax tillbaka , okej ? 
Allt kommer att bli bra . Mamma ska ta hand om dig . 
Min älskling . 
Du luktar som du igen . 
Vem skulle jag annars lukta som ? 
Det här kan brännas lite . Men det kommer att värma upp dig . 
Jag har saknat dig . 
Jag har saknat dig också . 
Åh , nej . Varmvattnet är slut . 
Jag ska koka mer . 
Gå inte . 
Mamma . Jag är kall . 
Mamma ? 
Var är du ? - Var är du ? 
Var ... - Jag är här . 
Vad är det som är fel ? 
Var är hon ? 
Vem ? 
TsUP , det här är Stationen . Uppfattar ni ? 
Hör ni mig ? 
Jag har förlorat tid . Jag har förlorat timmar . 
Jag tror att min syrenivå är låg . Jag svimmade i ... 
Återstående livsuppehållande , sex timmar och 45 minuter . 
Major Lysenko . 
Befälhavare Caldera . 
Du gör mig märkligt bättre till mods . 
Du säger alltid det , men jag vet aldrig om det är sant . 
Jag har utrustning här som omgående måste skickas med sök och räddning för Sojuz 1 . 
Det är osäkert om det blir nån sök och räddning för Sojuz 1 . 
Varför ? 
Vi får inga livstecken . 
Nu åker vi . 
Okej . Gör det . 
Det kommer att gå . 
Lugnt och fint . Lugnt och fi ... Ja . 
Jag vet inte om ni kan höra mig härifrån . Det här är Stationen . Batteri två är överfört till Sojuz . 
Det har tagit cirka 55 minuter att byta ett batteri . 
Jag har fyra kvar . 
Och sen 90 minuters avdockningsprocedur . 
Kan nån höra mig ? 
Det här är Stationen . 
Jag är mörkrädd . 
Det finns väl andra raketer ? 
Alla de där galna miljardärerna . StarCosm . Visst ? 
Även om StarCosm arbetar frenetiskt , kan de aldrig skjuta upp på knappt en dag . Och hon har inte en dag . Hon har några timmar . 
Det måste finnas ett sätt att få hem henne . Det måste vara möjligt . 
De hann inte skicka utträdesparametrarna i tid . 
Vad är en utträdesparameter ? 
Det betyder att även om hon lagar kapseln , måste hon kalkylera sitt eget återinträde . 
Det här är väldigt farligt . 
Men hon är tränad för det här . 
Jag menar , du tränade henne i fyra år . 
Åh , för guds skull , gråt inte . 
Sitt för fan inte där och gråt . 
Alice ... Är du klar ? 
Jag måste bara prata med de andra innan de åker . 
Är hon död ? 
Hon har inte mycket tid . 
Hon är väl inte död förrän vi vet att hon är död ? 
Jag älskar dig , gumman . 
Hej , älskling . Hej , Magnus . Jag tänkte att jag kunde spela in nåt eftersom jag inte kan prata med er . 
Okej , så jag måste fixa allt det här så att jag kan komma hem . 
Så konstigt att det liksom känns skönt att höra en röst även om det bara är min egen . 
Det här är det tredje . 
Jag måste skynda mig . 
... är det tredje . Jag måste skynda mig . 
Du måste sluta andas . 
Sluta andas , Jo . 
Stanna i Destiny . 
Paul ? 
Vad i helvete gör StarCosm ? 
Vi pratar med Alyanna . De försöker verkligen , men , Henry , hon hinner dö innan dess . Det är en svindlande summa pengar för att få hem två döda kroppar och lite experimentutrustning . 
Lite experimentutrustning , Michaela ? Det är oerhört betydelsefullt forskningsmaterial . Inte bara för vår teoretiska förståelse av universum , utan även för cirka tusen olika praktiska tillämpningar som kan göra en fundamental skillnad för livet på den här planeten . 
Vetenskapen kan inte trumfa människorna , Henry . 
Det här är TsUP . 
Hej . Uppfattat klart och tydligt . 
Nån chans för ett samtal med min familj i dag ? 
Stationen , det här är TsUP . 
Det här är en inspelning . 
Vi har S-frekvensavbrott och kan inte höra dig . 
- Öppna alla frekvenser för lokalsändning . 
Vi försöker ladda upp dina utträdesparametrar . RPL begär att du räddar CAL:s datakärna . 
Återställ full elförsörjning till Sojuz 1 . Initiera avdockning snarast . 
Du har cirka två timmar och 30 minuter av livsuppehållande från och med kl 9 : 38 den 15 / 10 . 
Kom igen . 
Stationen , det här är TsUP . Det här är en inspelning . 
- Öppnade ni kretsar ett och fyra ? 
- Ja . Det finns inget nära henne , inte från oss . 
Vi placerar inte satelliter i närheten av ISS . 
Oss emellan , amerikanska flygvapnet har flyttbara satelliter . 
Jag har bett dem placera dem högre . Vi vet det , Henry , men att flytta dem närmare hjälper oss inte att nå henne . 
Om skadorna är för betydande , kan hon kanske inte höra längre . 
Befälhavare Caldera , ni har ett samtal från Skagerrak marinobservatorium . 
Åh , jisses . 
Skagerrak ? 
Se inte på mig så . 
Jag tänker inte förlora varken CAL eller henne . Så blir det inte . 
Stationen , TsUP . Det här är en inspelning . 
Vi har S-frekvensfel och kan inte höra dig . 
Har du hört från din syster ? 
Jag tror att du vet att hon är död . 
Har du hört från din bror ? 
Inte på många år . 
Tack och lov . 
... inväntar besked om vad som hänt astronauten som är kvar på ISS ... SS BERNICE 12 SJÖMIL UTANFÖR KALIFORNIEN ... nu bokstavligen den ensammaste personen i universum . 
Med mig har jag pensionerade astronauten Bud Caldera . 
Befälhavaren , vad händer när strukturen på ISS skadas på det viset ? Det skulle leda till en " depress " , tryckförlust i de olika modulerna på ISS . Det är i stort sett det allvarligaste som kan hända . 
Beskriv vad som troligen pågår där uppe med den kvarvarande astronauten . 
Det följer ett regelverk . 
Vi har blädderböcker med checklistor , och vi går igenom i stort sett varje scenario under utbildningen . 
Så även om det är en ovanlig situation , arbetar de enligt en plan . 
Men ni har erfarenhet av vad som kan hända om nåt går snett där uppe . 
Visst . 
Det måste locka fram en del minnen . 
Nej , jag söker inte efter ... Jag ödslar inte min tid på minnen . 
Men ni har erfarenhet av hur det är att föra hem kroppar . 
Det är ingen fråga . Det är en observation . 
Kan ni kanske bara berätta lite om hur ni tror att de känner just nu ? 
Ja , och varför i helvete skulle jag det ? 
Och säg mig vad " lite " är . 
Jag får inte betalt för att använda min satans fantasi . 
Henry Caldera , stort tack . 
Jag heter Bud ! Bud Caldera , för guds skull . 
Helvete . 
TsUP , det här är Stationen , kom . 
Elförsörjningen är fullt återställd på Sojuz 1 . 
- Stationen , det här är TsUP . 
- Det här är Stationen , kom . 
Det här är en inspelning . 
Du har cirka 98 minuter livsuppehållande från och med kl 10 : 48 . Avdockningstid är minst 90 minuter . 
RPL begär att du hämtar CAL:s datakärna . Du skojar . 
Vi försöker ladda upp dina utträdesparametrar . 
Jag kan inte vänta . 
Kom igen . Kom igen , kom igen , kom igen , kom igen . 
Vad i ... " Syre : 19 % . " 
Jag måste iväg . 
I blindo . 
Initierar avdockningsprocedur , Sojuz 1 . 
" Mata in utträdesparametrar . " 
Jag använder gårdagens siffror , för det är allt jag har . 
" Utträdesparametrar förlegade . " 
Ja , jag vet , men du måste samarbeta . 
Åh , kom igen . 
Kom igen , kom igen . Snälla , kom igen . 
" Avdockning initierad . 
Nittio minuter till uppskjutning . " 
Stationen , det här är TsUP . 
Det här är en inspelning . 
Vi har S-frekvensfel och kan inte höra dig . 
Var snäll och öppna alla frekvenser för lokal sändning . 
Vi försöker ladda upp utträdesparametrar . 
Pappa , vad är utträdesparametrar ? 
Som jag förstår det , är det platsen i utkanten av jorden som man måste pricka in om man vill komma hem . 
Vet mamma vad de är ? 
Jag vet inte . 
Det vet hon säkert . 
Hon är väldigt smart . 
- Håll käften . Vi har S-frekvensfel och kan inte höra dig . 
Var snäll och beräkna dina egna utträdesparametrar . Det har jag gjort . 
RPL begär att du räddar CAL:s datakärna . - Försätt dig inte i fara . - Åh , för helvete . 
Hej , Magnus . 
Jag ska mata in utträdesparametrarna . Mina egna beräkningar . 
Låt oss bara hoppas att de tar mig hem . 
Fyrtioett ... Magnus , jag känner dig . Och du vet varför jag måste göra det här . 
Och jag är så tacksam för din kärlek och din tillit . 
Jag vet att det inte har varit lätt . Du har offrat mycket ... Jag är ledsen att jag jag lämnade dig ensam med allt det här ... 
Jag älskar dig . 
Du är mitt allt . 
Och jag ville ... Jag ville göra dig stolt . 
Dig . 
Och jag ville visa dig att ... Även om jag inte är här så finns jag alltid hos dig och pappa . 
Jag tror inte att du förstår hur mycket jag ... Jag ville bara finnas där och se dig växa upp och gå på gymnasiet och ha din första pojkvän och och sen gå ut och dansa med dig när du blir vuxen och bara ... 
Oavsett vad som händer , så är mina ögon alltid på dig . 
Och mitt hjärta slår med dig , älskling . 
Jag älskar dig så mycket , mer än du nånsin kan ana . 
Okej . Så , jag har bara 12 minuter kvar , och jag måste liksom ... Jag hoppas bara att jag har räknat rätt . 
" Bultfel " ? 
Vad ? Vad fan ? 
Armbultarna är i funktion . Kan inte vara uppgifterna . 
" I händelse av bultsystemfel , ska bultar laddas och avfyras från ISS:s ingångsbrygga på andra sidan luckan . Kräver två besättningsmedlemmar . " Helvete . 
Kom igen . Kom igen , snälla . 
Fyrtioett , 40 , 39 , 38 , 37 , 36 , 35 , 34 ... Nån trianguleringsinformation ? Inget . Fortfarande inget . 
... 30 , 29 , 28 , 27 , 26 , 25 , 24 , 23 , 22 , 21 , 20 , 19 , 18 , 17 , 16 , 15 14 , 13 , 12 , 11 , tio , nio , åtta , sju , sex , fem , fyra , tre , två , ett . Lyssna . 
Slut era ögon . 
När namnen på dem som somnat in koms ihåg i böner , vad kan vara mer välgörande för dem än det här ? 
Vi som lever tror att de döda inte har berövats sin existens , utan lever med Gud . 
Såsom vi ber för våra bröder och systrar som med tillförsikt och hopp reser , ber vi för dem som har lämnat denna värld . 
Jo , det här är TsUP . 
Uppfattar du ? 
Lossad från ISS . 
Tre timmar och 20 minuter till återinträde ... Tror jag . 
Jag tänkte att du kanske inte ville vara ensam . 
Jag är ganska tillfreds med att vara ensam . 
Så , hur mycket tar ni för en tur-och returresa på Sojuz numera ? 
Sjuttiofem miljoner , upp och tillbaka ? 
Det lider mot sitt slut . 
Såvida ni inte börjar skicka turister . Turister ? 
Åh , snälla . 
Skål . 
För Jo och Paul . 
Avfyrar om fem , fyra , tre , två , en . 
ISS skapades inte för att hållas i drift längre än 20 år . Den har hållits i drift i nästan 30 . 
Och den är full av hål . 
Din egen president säger högst sju år till . 
Min egen president har fel . Jag jobbar på min egen president . 
Vi kommer att dra oss ur programmet . 
Bara överge saker för att nåt gick snett , för att nån dör ? 
NASA övergav månen efter Apollo 18 . 
Så det är vad det här handlar om ? 
Du vet vad jag har sysslat med i alla dessa år . 
För mig handlar det kanske om det . 
För Roskosmos handlar det om att utnyttja ett naturligt avslut . 
Är du inte minsta nyfiken på sjukdomen på vilken du är en expert ? 
Det skedde en dödlig olycka efter åratal av varningar om rymdskrot . 
Det här kommer att hända igen , Henry . 
Och det finns en stor mängd svar som vi aldrig kommer att få . 
Jag håller med . Vi utnämner ISS till en internationell grav , och överlåter rymden åt människorna med pengar . 
Sojuz 1 , det här är TsUP . Hör du mig ? 
TsUP , det här är Sojuz 1 i återinträde . Uppfattar ni ? 
Det här är Sojuz 1 , kom . Snälla . BALLISTISK LANDNING KORRIGERA KURS OMEDELBART 
Sojuz 1 har återinträtt i jordens atmosfär . Hon svarar inte . Den inträder ballistiskt . 
- Var slår hon ner ? - Varsomhelst inom 300 kilometer . 
Ta fram era amatörradior och hitta henne . Vi måste ta reda på var i helvete hon är . 
- Det är en nål i en höstack . 
- Kan du inte ringa NORAD ? Ring din jävla kille i Egypten . 
Roskosmos markkontroll , Sojuz 1 här . Hör ni mig ? Roskosmos markkontroll , Sojuz 1 här . Hör ni mig ? 
Sojuz 1 ... Sojuz 1 , det här är TsUP . Hör du mig ? 
Sojuz 1 , det här är TsUP . - Vi hör inte ... - Fan . - Öppna alla VHF-frekvenser . 
Sojuz 1 , det här är TsUP . Upprepar . Öppna alla VHF-frekvenser . 
Det är en ... Jag försöker ! Jag försöker ! 
Sojuz 1 , vi hör dig . 
Du har avvikit 6,5 grader från optimal kurs , du måste korrigera . 
Jag är i ballistiskt inflygningsläge . Jag kan inte . 
Fråga om hon hämtade datakärnan . 
- Åh , Henry , för guds skull . 
- Fråga henne . Har du CAL:s datakärna ? Ja . 
Har ni henne ? Var är hon ? Du flyger in i väldigt brant vinkel . 
Du når snart 8G . 
Förstått . 
Jo , du försvinner . 
Det lär ta tid att hitta dig . Lycka till . 
Hej . Vet du vad ? 
Vad ? 
Den är märkt med RPL-blixtar . Den ska med sök och räddningshelikopter 1 . 
- Sätt fart nu , för helvete . - Ska bli . 
Hon har superkort tid . Det blir väldigt svårt att hitta henne . 
Gör inte så här mot mig , Frederic . Jag har just lugnat min dotter . 
Vi flyger åt nordost men ser inget från helikoptrarna . 
Helikopter 5 , kolla sydösterut ovanför berget . 
Helikopter 2 , nordväst 22 grader . 
Fortfarande inget , Team 1 . 
Mamma ! 
Det är min älskling . 
Sätt ner mig . Sätt ner mig . Det är min älskling . 
Mamma ! 
Jag älskar dig . 
Jag älskar dig så mycket . 
Är du okej ? 
Jag är så ... Jag är så glad över att vara här . 
Jag älskar er så mycket . 
Jag älskar er så mycket . 
Jag ... Välkommen tillbaka . 
Tack . 
Ge mig den , tack . 
Öppna kapseln . 
Behållarna borde vara iordninggjorda . 
Det här är mitt skötebarn . 
Ge mig iPaden . 
Ge mig lite utrymme . ANSLUTER 
Är det Wendys pappa ? Du behöver inte titta , älskling . Titta inte . 
Så , hur är det ? 
Jag vet inte . 
Åh , du ser fantastisk ut . 
Jag är tillbaka . Jag tog mig tillbaka . Ja . 
- Hej . Jo , jag ... 
- Kom . Nu går vi . 
Sätt fart , hörni . 
Jag är strax tillbaka , älskling . 
- Jag är tillbaka nu . - Hon är hemma . 
Vi kör dig direkt till Star City . 
Ursäkta . 
Lägg undan kamerajäveln . 
Herrejävlar . Den är där . 
För helvete . 
Den kan inte vara där . 
Hur säger man " heureka ! " på ryska ? 
Mamma ? 
Är du okej ? 
Vad ? 
Man glömmer hur jorden luktar . 
Var är hon ? Vem ? 
Var är min älskling ? Alice ! 
- Vad ? - Var är hon ? 
- Vem ? 
- Du . 
Jag vet inte vad du menar . 
Såg du inte dig själv ? 
- I spegeln ? - Nej ! Här . Mamma , jag såg inget . 
Klä på dig . 
Mamma ! 
Gör dig klar . 
Kom , vi måste iväg ! 
Det är för kallt . Hon fryser ihjäl . Vi måste hitta henne . 
Vem ? 
Den andra du . 
