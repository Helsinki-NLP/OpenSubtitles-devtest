Hej , det är Kyra ! Välkommen till min kanal . 
Glöm inte att gilla och prenumerera för jag lägger upp nya rese - och matvideor varje dag , och ni vill inte missa dem . 
Jag ser fram emot vårt nästa resmål , Philadelphia ! 
- Gör du det också ? - Jag gillar att vara med dig . Ifall det inte var uppenbart . 
- Jag älskar dig . 
- Detsamma . - Vad vill du äta ? - Jösses ! 
Allt . Matscenen i Philly är grym . 
Vi ska testa trendiga ställen och streetfood . - All mat är god , oavsett budget . - New York blir svårslaget . 
Ja , men jag ser fram emot Philly-kringlan . Och sorbet givetvis . Jag kan inte sluta tänka på Philly cheesesteak . 
- Nu gör du mig hungrig . 
- Mig också . 
Jag taggar alla ställen på Insta . @ KruisingWithKyra . Kruising med " K " . Följ mig där om ni vill ha alla rekommendationer . 
Philly är så vackert . 
Min mormor och morfar träffades här . Vem vet , Teddy kanske friar till mig här . - Kyra ! Seriöst ? - Våra följare älskar det . 
Nej , dina följare gör det . 
Varje gång du nämner förlovning får jag skit . 
" Teddy vet inte vad han har . " " Teddy , sätt en ring på fingret . " 
" Varför är hon med honom ? Han är medel . " - Det är inte roligt . 
- Förlåt . Jag försöker bara bygga nåt åt oss båda . 
Jag bad dig att radera klippet från Central Park . 
- Jag såg ut som en idiot . - Nej . 
Det är det enda klippet jag har på oss två . 
Jag tar bort det . 
Vad är poängen ? Det har redan 50 000 visningar . 
Börja om . 
Hej , det är Kyra . Välkommen till min kanal . 
Glöm inte att gilla och prenumerera . Jag laddar upp nya rese - och matvideor varje dag . 
Jag ser fram emot vårt nästa resmål , Philadelphia ! 
- Hej . Proviant . 
- Är du galen ? 
Det ösregnar ! 
- Jag mår bra . Hur mår du ? - Förlåt mig . 
- Är du galen ? 
Det ösregnar . 
- Väldigt gulligt . Skulle inte du träffa snubben som erkände bilbombningen ? 
Logan Barlowe . Vägen till Frackville är översvämmad . - Jag fick boka om . - Ost , kex , vin och ljus ? 
- Ja , sånt jag hade hemma . 
- Sånt du hade hemma ? 
Jag måste säga att jag gillar det här . 
Du behöver lite saker på grund av stormen . 
Du organiserade svensexan åt din exfrus nye man . Hur gick det ? 
- Du behöver inte göra så . 
- Vad då ? Du gör det konstigt med dina ord . 
- Mina ord gör det konstigt ? - Ja , dina ord . 
- Menar du mina fakta ? 
- Mike är min partner och vi hade kul . 
- Toppen . Hade Nikki kul ? 
- Jag vet inte . 
Det ligger en kropp på baren . - Jag är här . 
Har festpatrullen varit här ? 
Ja , du vet , vår ursprungliga plan spolades bort . 
Du borde städa innan Braun får veta nåt . 
Han gav mig sitt godkännande . Han till och med bidrog med champagne . 
Var han snäll för en gångs skull ? 
Vilken tur att du sov här , jag kunde knappt ta mig in . 
Vi kanske var lite väl entusiastiska . 
På en skala från ett till Chocolate City ? 
- Jag har inte frågat om din fest . 
- Är det reglerna ? 
Ja , möhippor är heliga . 
Då säger jag inte vad jag och Jay gjorde . 
- Helt okej . 
- Vidrigt . 
- Kaffe ? 
- Kaffe . Vakna , Helen ! 
God morgon , kriminalinspektör Sherman . 
- Jösses ! 
- Hej . - Du vet väl att vi äter på den . 
- Hjälp ! Jag behöver hjälp ! Jag vill anmäla en försvunnen person . 
- God morgon , solstråle . 
- Sluta . Filma mig inte utan smink . 
- Du är perfekt som du är . 
Vart för våra äventyr oss idag ? 
Ni ser så glada ut . Hur länge har ni varit ihop ? 
Två år . 
Vi träffades på en fest i college . Vi pratade om platser vi ville besöka , musik , livet . Hon är lätt att prata med . Kyra får alla att känna sig speciella . 
- Och ni bor i en skåpbil ? 
- Ja . 
Efter examen hade Kyra redan många följare . Hon la upp videor på YouTube och TikTok . Matrecensioner och resor . 
Vi bestämde oss för att renovera skåpbilen och resa . 
Planen var inte att bo i en skåpbil men jag skulle bo i en grop med henne . 
- När kom ni till Philadelphia ? 
- För tre dagar sen . När jag kom tillbaka imorse var hon borta . 
Och skåpbilen var borta . 
Det går inte ihop . 
Teddy , finns det en chans att Kyra bara behövde en paus ? 
- Ni kanske bråkade ? 
- Nej . Är du säker ? 
Det är tufft att bo så trångt . 
Nej , vi älskar varandra . 
Jag vet att nåt har hänt henne . 
Känner Kyra nån i Philly som hon kanske hälsar på ? 
Nej , och hon svarar alltid när jag ringer . 
- Har du kontaktat hennes föräldrar ? 
- De är döda . Hennes mamma dog i cancer , hennes pappa kort därpå . 
- Kyra sa av brustet hjärta . 
- Det låter tungt . Hon har ett hål i hjärtat där hennes föräldrar brukade vara . 
Hon vill ha många följare för att fylla det tomrummet . 
- Jag försökte . 
- Jag lovar att göra allt vi kan . 
Sen hennes föräldrar dog avskyr hon att vara ensam . 
Det skrämmer henne . Hon skulle aldrig sticka sin väg . 
Jag vet att nåt hemskt har hänt . 
Följ med mig , så ska du få torra kläder . 
I den här stormen tar jag inga risker . 
Jag efterlyser Kyra . 
FÖRSVUNNEN - Försvunnen flicka . Jag måste gå . 
- Det är orkan där ute . 
Jag vet , men det är mitt jobb . 
Det är vad jag gör , så jag måste göra det . 
Jag kommer tillbaka senare och tittar till dig . 
Jösses , vad män är korkade . 
Glömde du manteln , supersnuten ? 
Det var roligt . 
- Duschar du med kläderna på ? 
- Jag såg Kyras efterlysning . 
Hennes pojkvän anmälde henne försvunnen imorse . 
Är du på Waynes motell ? Flott . 
Festen slutade visst sent . 
Nej , han tittade bara förbi . 
- Med proviant . 
- Proviant . Kan du hämta mig ? 
Min bil är under tre meter vatten . Omöjligt . Guvernören utlyste undantagstillstånd . 
Floden är översvämmad . 
Hela byggnaden är avspärrad . 
Vilken idiot stänger ner polisens högkvarter ? 
- Låt mig gissa . 
Braun . - Jag vet inte . 
Men det är galet där ute . Jag vet inte hur vi ska hitta Kyra . 
Okej . 
Vad gör vi nu ? 
- Är du okej ? 
Kyra De la Cruz , 22 år . Reseinfluencer . 
Sågs senast imorse nära centrum av sin pojkvän , Teddy Williams . Jag söker på trafikkameror efter deras skåpbil men det är dålig sikt i det här vädret . 
- Efterlysningen gav inget . 
- Eller hennes mobil . Den är avstängd eller stulen . 
Gräv i Kyras sociala medier efter ledtrådar , platser , fanatiska fans . 
- Kan jag hjälpa till ? 
- Helen ? - Ja , chefen . Kan du ta med konstapel Hardbody nånstans som inte är här ? 
- Javisst . 
- Tack . Mitt riktiga namn är Jack . 
Eller Jackson . Konstapel Hardbody är mitt scennamn . 
- Det förvirrar mig också . 
- Helen ! 
Förlåt . 
- Kom igen , Jack . 
Vi säger till när nedstängningen är hävd . 
Jag kan inte ta honom på allvar i den lilla västen . 
- Jösses ! 
- Vad händer ? 
Teddy bad följarna på Insta om hjälp att hitta Kyra . 
Tipsen strömmar in . 
Be alla lediga poliser om hjälp . Det är goda nyheter . 
- Konstapel Hotpants också ? 
- Någon vet något . 
Jag vill ha en rapport på mitt kontor om en timme . 
- Har nån sett Jay ? 
- Ja , Waynes motell . 
En tjej är i knipa och jag är fast här och spelar kort . 
Sju kort . 
Du kastar och drar ett kort varje gång . 
Man samlar fyrtal och tretal , antingen i samma valör eller färg . 
- Då har man gin . Förstått ? - Uppfattat . 
- Hej . - Jag är fortfarande fast på motellet 
- Ska jag simma till jobbet ? 
- Han bör vänta ut det . 
Hon har rätt , Jay . 
- Vi jobbar på det . 
Jag hörde att du flyttade möhippan till MPU . 
- Vad gjorde du och Mike ? 
- Det säger jag inte . Han sa att jag inte fick säga nåt . Något om en bro-kod . 
Herregud ! Ni och er bromans . 
Lova att inte göra nåt galet . 
Jag märkte att du inte lovade att inte göra något galet . - Inte det ? 
- Jason Grant vill inte vara bunden . 
- Eller så gör han det . Vet inte än . 
- Väldigt lustigt . 
Om du hade din laptop hade vi kunnat hjälpa tjejen . - Jag säger bara . 
- Min laptop . Flytta på foten . 
Du tar Supersnut-grejen bokstavligt . Det är lustigt . 
Den var i bakluckan . Snyggt . 
Då kör vi . 
Starta den , så ska vi se om vi kan hjälpa Kyra . 
Den behöver laddas . 
Den jäveln . 
Sen såg jag att Kyra twittrade motsatsen bara en månad tidigare . 
Jag vet inte , men det verkade misstänkt . 
Rome , det är toppen . 
Vi har dina kontaktuppgifter och hör av oss . 
- Nik ! 
- Vad har du hittat ? 
Det här är Rome Carter-Lee . Välkomna till " True Crime " med Rome . 
En liten uppdatering om Kyra De la Cruz . 
Han är från Philly och har ringt in tre gånger . 
Är han ett fanatiskt fan ? Han har en brottsblogg på TikTok och verkar äkta . - Dömd för trakasserier och stalking . 
- I vilket sammanhang ? 
Offret var en lokal influencer som ansökte om kontaktförbud . 
Vi tog bort hans sista objekt . 
Han kanske fick ett nytt i Kyra ? 
Han la upp en video om henne . Han säger att hon fejkar sitt eget försvinnande . 
- Och kritiserar Teddy . 
- Arg , svartsjuk och fixerad . 
Frågan är bara om det är mycket snack och lite verkstad . 
Kemi får kolla upp det nu . Den här mannen är farlig . 
- Rör den inte ! 
- Vad är det ? En hybridiseringsinkubator . 
Hybrid ... inkubator . 
Du är så smart . 
Rör inte den heller ! 
- Du ... 
- Jackson . 
Jag vet att du sitter fast här också , men det här är mitt jobb . Det är min arbetsplats . 
Jag är ny och jobbar hårt för att få alla att gilla mig lite . 
Varför skulle de inte gilla dig mycket ? 
Sitt där borta tills stormen är över och låt mig jobba . 
- Gillar du musikaler ? 
- Gillar dem ? Jag älskar dem . 
Jag spelade Fiyero . 
Så du är ... Jag trodde att du var ... Min lillebror är gay . 
Heterokillar gillar också musikaler . 
- Var min kyss så hemsk ? 
- Kysstes vi ? - Vi kysstes . 
Vi kysstes . 
- Den var het . 
- Jag dricker aldrig champagne igen . 
Ta den här ! Och gör en lista på alla svåra saker som ... 
Uppför dig ! Annars låser jag in dig i förhörsrummet . 
Det vore inte så illa . 
Ett batteri , en växelriktare . 
- Fantastiskt . 
- Är du säker på att det funkar ? 
- Bara den inte läcker vätgas . 
Jag kanske borde flytta ljuset . 
Nu jobbar vi på att hitta flickan . 
- Kan jag göra något ? 
- Den är blöt . 
- Du har rätt . Det är bara en ledare . 
Det är okej . 
Det funkade . 
Romes teorier om Kyras fall är logiska . 
Antalet följare har fördubblats . Men det har hans också . 
Han utnyttjar och kränker henne på samma gång . 
Sen hittade jag det här . En taggad bild på Instagram . 
Rome träffade Kyra för tre år sen på TrendingCon . - En konferens för influencers . 
- Han glömde nämna det . 
Enligt kommentarerna började de gräla . 
Och när Kyra besöker hans hemstad försvinner hon . - Vi verkar ha oss en misstänkt . - Ja , det har vi . 
Det är Jay . 
- Hej ! Det är fler ljus än på din senaste födelsedagstårta . Jätteroligt . Strömmen gick , men vi är tillbaka . 
Nåt nytt ? Rome Carter-Lee . Besatt av brott och har Kyra-problem . 
- Jag kollar honom . - Bra . 
Vi har en dömd stalker . Hon kanske gick rakt in i en fälla . 
Kan du förklara varför du är på ett foto med en försvunnen flicka ? Som du nu utnyttjar för fler visningar ? 
Jag träffade hundratals personer . 
Hade jag kommit ihåg det fotot , så hade jag använt det . Vi bryr oss inte om dina inlägg , utan om dina tidigare domar . 
Minns du Emily Beck ? 
Den subban försökte få mig blockerad . 
" Subban " ? Din mamma måste vara stolt . 
- Det här är illa . 
- Vad då ? 
Våra kollegor kan se att du beställde boken , " Sanering av brottsplats " . 
Behöver du sanera , Rome ? 
Jag söker på morbida saker för min TikTok-sida . 
- Men jag skadade inte Kyra . 
- Det vet man aldrig . 
Jag är inte er kille . Det handlar alltid om tre saker . Slumpen , brott , olycka . 
Och det faktum att er försvunna tjej precis la upp en ny video , så gissar jag att det är den första . 
Kan ni komma hit en stund ? 
Rome hade rätt . 
En ny YouTube-video kom precis upp . 
Hon måste ha förinspelat den och schemalagt den idag . 
Det är rätt vanligt bland vloggare . 
Hejsan ! Jag börjar med att säga att ni inte ska oroa er för mig . 
Det ser ut som om jag har gråtit , eftersom jag har det . 
Teddy och jag bråkade , och jag behöver bara lite egentid . 
Teddy sa att de inte bråkade . 
Han sa även att de sågs imorse , och sist solen sken var igår . - Den spelades in då . 
- Så han ljög om när hon försvann ? 
Att anmäla henne försvunnen är ingen dålig plan om man vill lura polisen . 
Drömprinsen verkar ha en del att förklara . 
Kommentarerna fullkomligt exploderar . 
" Teddy , hur kunde du ? " " Vad gjorde du med Kyra ? " 
- Till och med dödshot . 
- Internet skiftar snabbt . 
Be Helen DNA-testa Teddys blöta kläder . 
Jag tror att vår kille har lurat oss . 
Teddy och jag bråkade . 
Jag vet att det ser illa ut . 
Det är illa att du sa att ni sågs imorse . 
Att ljuga om ett bråk är väldigt illa . - Var är hon ? - Jag vet inte . 
- Är hon skadad ? 
Lever hon ? 
- Jag vet inte ! - Vi bråkade igår . 
- Om vad då ? 
Hon ville lägga upp ett inlägg om förlovningsringar och jag kände mig pressad . 
Det är nog läge för dig att skaffa en advokat . 
Du lyssnar inte . Jag älskar henne . 
Jag har inte gjort nåt . 
Han är orolig . 
Frågan är varför . 
Hashtaggen " Hitta Kyra " trendar . 
Alla vill ha en del av dramat . 
De är bara sensationslystna . 
Vi måste fastställa när hon försvann . 
Jag har kartlagt hennes sista timmar via hennes digitala fotavtryck . 
Kl . 10.00 på söndag lägger Kyra upp deras ankomst i Philly på Instagram . 
Kl . 12.13 lägger hon upp på TikTok att hon äter en kringla vid Liberty Bell . 
Kl . 14.41 tar ett fan en bild med dem båda på John ' s Water Ice . 
Kl . 19.00 twittrar Kyra från middagen på Locus på Rittenhouse Square . 
Och till sist , kl. 08.00 på måndagen på Kyras Instagram-story : " Vaknar i Philly " . Och de ser ut som två glada campare . 
Så de bråkade efter det . 
Minns du den nya YouTube-videon som hon la upp ? 
Vi vet höjden på lyktstolpen i bakgrunden . 
Via skuggans längd kan jag räkna ut att videon spelades in cirka 11.00 . 
- Du är grym . - Tack . Det betyder att de grälade mellan kl. 08.00 och 11.00 igår morse . 
Ja , och det finns ingen annan onlineaktivitet förrän kl. 17.32 då hon lägger upp en BeReal från en bar i Kensington . 
- BeReal ? 
Den skickar ut notiser som ber användaren att lägga upp ett foto inom två minuter . Poängen är att det är spontant . 
- Man såg att hon hade gråtit . 
- Och sen är hon borta . Det betyder att den senast kända platsen var Kensington . 
Nåt mer ? Det är en chansning , men om vi kan se hennes opublicerade videor ... 
Vi letar efter en opublicerad video som visar vart Kyra gick efter sitt inlägg igår kl. 17.30 . 
- Jag hackar molnet nu . 
- Vi kollade upp Rome Carter-Lee . 
Förutom att han verkar tro att Kyras försvinnande är hans stora genombrott som fåtöljdetektiv visar hans mobildata att han inte har lämnat sin mammas källare på en månad . 
Det betyder att Teddy är vår huvudmisstänkte . 
Jag har dåliga nyheter , inga schemalagda uppladdningar . 
Om videokameran har automatisk backup kan jag komma åt originalet . 
- Tillstånd att hacka ? 
Kom igen , vi behöver ett genombrott . 
Toppen , jag uppskattar det . Tack så mycket . En trafikpolis i Camden County såg efterlysningen . 
Han stoppade Kyra och Teddys skåpbil förra månaden . Ett bakljus var trasigt . 
Han försökte förhöra henne separat , men hon vägrade . - Misstänkte han misshandel ? 
- Han lät dem åka . Provsvaren på Teddy Williams kläder kom . 
- Jag fann en blodfläck på skjortan . - Hans eget ? 
Det är DNA från en kvinna . 
Vi har bilderna från kroppskameran på polisen som stoppade er . 
När en person tar hårt i sitt offer lämnar det såna här märken . 
- Tror du att jag gjorde det ? 
- Japp . Kyra föll under en fotvandring . 
Vi har videobevis . Jag skulle inte ... 
Du ljög om när ni såg sist och om ert gräl . 
Jag var rädd att ni inte skulle tro mig och tänka att hon dumpade mig . 
Hur förklarar du kvinnoblodet på tröjan du bar imorse ? 
Det är från fotvandringen . 
Vi ödslar tid när ni borde leta efter Kyra . 
Teddy ! Finns det någon där ? 
Hjälp ! Är det nån där ? 
Hjälp ! 
- Ja ? 
- Hej . Wayne hackade Kyras molnserver och fann en video från kl. 20.30 igår kväll . 
Trots alla tokigheter kunde jag inte komma hela vägen till Philly utan att äta en cheesesteak i ett av stans äldsta ställen . 
De gör sin variant av klassikern , så den är lite dyr men om jag ska äta mina känslor är jag på rätt spår . 
Är det koriander och fänkål ? 
Jag känner ingen ostsmak alls . 
- Är det taleggio ? 
- Stackars tjej . 
Jag ville bara att en sak skulle gå rätt idag , så jag unnade mig den här dumma , dyra mackan som suger . 
Ännu en gång tar en kock nåt vi älskar och försämrar det . Det här stället är inte värt pengarna . 
Vad fan sa du ? Spelar du in nu ? 
Stäng av kameran . Stäng av den ! 
- Du gör mig illa ! - Vem sjutton är det ? Identifiera honom . 
Så fort du kan . 
En helikopter ? 
Jag vet att du vill vara snäll , men det är onödigt . Jag mår bra . 
Ja . Vi vill vara diskreta och en helikopter är inte diskret . 
Jag måste gå . Hej då . 
Ville din mystiske man skicka en helikopter ? 
Vem är han ? Hon drack fyra tequilashots igår utan att säga nåt . 
Ni får träffa honom på bröllopet . 
Om han slutar att försöka rädda mig . Det är bäst för honom . 
Då ska vi se ... 
Kyras angripare är Nico Falcone från Falcone ' s Original . 
Stället öppnades av deras farmor Rose på 1930-talet . Det sägs att bröderna Olivieri uppfann cheesesteak men Rose fulländade den . 
Jag älskade deras " whiz wit " . Jag har inte varit där sen de ändrade familjereceptet . 
Du är inte den enda . 
Då ska vi se . 
Titta på det här . 
De ligger efter med hyran . 
Och det är inte allt . 
De har inte betalat elen på flera månader . 
Nico växte upp i Toscana . 
När hans farbror dog tog han över restaurangen och hade med sig några konstiga idéer . 
Wagyu-cheesesteak är en dummare än dum idé . 
- Det låter så . - Jösses . 
Han har maxat sina kreditkort och kan inte betala av ett lån . 
- Och han är tidigare straffad . 
- Innehav och grov misshandel . 
Så problem med ilska och droger och nära att förlora familjebolaget . 
Och in kommer Kyra och sätter en sista spik i kistan . 
Om stormen inte låter oss gå till Nico , så får Nico komma till oss . - Ja . 
Kom igen . - Hallå ? 
Känner jag er ? - Kriminalkommissarie Batista . 
- Jag har inte tid att prata . - Det är brådskande , mr Falcone . - Nej ! 
- Strömavbrott . 
Vi har äntligen en misstänkt och strömmen gick . 
Jag såg videon . Han är våldsam och tidigare straffad . 
Det är illa . Vi kan inte göra mer förrän stormen är över . 
Jag kan ta mig till Falcone ' s. Nej , staden är översvämmad . 
Stanna ... - La du på ? 
- Vad ska jag göra ? 
Någons barn är i trubbel . 
Ska jag bara sitta här ? Du gillar inte att följa direktiv . Påminn mig om vem som bär fotboja . 
Du eller jag ? Det är jag . Och till och med jag vet att ibland är det bara smartast att sitta ner , hålla tyst och vänta på rätt tillfälle . 
Vänta på rätt tillfälle ? 
Minns du flygresan från Kandahar ? 
Arton timmar på ett plan och oroa sig över Keith . Undra var han är utan att kunna göra nåt . 
Jag tänker inte sitta i det här motellrummet när någons barn är i trubbel . Jag gör det bara inte . 
Falcone ' s är 10 kvarter bort . 
Visst , vill du drunkna ? Varsågod . 
Hallå , någon ? Hjälp ! Någon ? 
Nej ! Hjälp ! 
Hjälp ! 
Teddy ! 
Det är bara tio kvarter bort . 
Hur fan tänkte du ? 
Du har ingen plan , ingen backup . 
Du vet inte vad du ger dig in på . 
Jay ? Jay ? 
- Herregud ! 
- Vad är det ? 
Han går till Falcone ' s. Jag har fått nog av honom . Slappna av . Det blir ... 
Vill du ha en proteinshake ? 
Tragiske Mike , vill hon ha protein , så fixar Big Mike det . 
Och knäpp skjortan . 
Vi letar efter en saknad person . 
- Vi har stängt . - Philadelphiapolisen . - Jag gillar inte dyra mackor . - Toppen , gå till en Micky D ' s. 
Jag letar efter en tjej som heter Kyra De la Cruz . 
- Vet du vem det är ? - Ingen aning . 
Hon kom in igår kväll och gjorde en liten video . - Du attackerade henne . 
- Är allt bra ? 
Det beror på vem man frågar . 
Hon dissade min mat , jag gjorde sönder hennes kamera . 
Det handlar inte om kameran . 
Hon är försvunnen . 
Misshandlar du alla dina kunder eller bara dem som klagar på maten ? Är hon försvunnen ? 
Tror du att jag ... Du har fått det om bakfoten , amico . 
- Har jag ? 
- Ja . Vad har hänt med din skåpbil ? 
- Jag vet inte vad du pratar om . 
- Vad heter du ? 
- Johnny . - Läget , Johnny ? 
Mår du bra ? 
- Ja . - Tar du droger , Johnny ? - Nej . 
- Varför skakar du och är så nervös ? 
- Jag mår bra . Vad är det med dig ? 
Du måste svara , jag är polis . 
Berätta vad det är . 
- Jag tänkte säga nåt . 
- Vad då ? Efter du slog sönder kameran bad jag henne radera videon . 
- Vad fan , Johnny ? Vad gjorde du ? 
- Hon har en miljon följare . Det sprider sig snabbt . 
Så jag följde efter henne . 
Följde du efter henne ? 
Vad hände sen ? Jag tappade besinningen . 
Jag var arg . Jag prejade henne och hon körde av vägen . 
- Vad fan , Johnny ? 
- Lämnade du henne där ? 
Det var en olycka . 
Jag borde ha stannat , men ville inte få problem . Vad kallar du det här ? Du kan ruinera oss . - Var hände det ? 
- Nånstans i Fishtown . 
- Vad händer ? 
- Kemi , gör mig en tjänst . Kolla alla trafikkameror från igår i Fishtown . 
- Kyra prejades av vägen . 
- Uppfattat . 
Nikki ! 
Restaurangen är stängd . 
Stanna här tills tjejen är i säkerhet . 
Och Wagyu-cheesesteak ? 
Vart ska jag , Kemi ? 
Vi har fortfarande ingen ström , så jag vet inte , Jason . 
- Vad har de gjort med henne ? - Lugna dig . Kemi är bäst . 
Förlåt att jag avbryter , men jag kör i blindo . 
- Vi jobbar på det . 
- Ni kan inte hitta henne . 
- Strömmen är tillbaka , Jay . - Utmärkt . Prisa gudarna ! 
Det här ser bra ut . 
- Fishtown är en labyrint . 
- Nu börjar det likna nåt . 
Öster om floden , nära motorvägen . 
Hon verkar ha voltat ner i floden . - Herregud . 
- Lyssna på mig . Jason och jag har en dotter i Kyras ålder . 
Han gör allt för att se till att hon är säker . - Vad gör du ? 
- Jason är jobbig . Men han är min partner . Om han går , går jag . Bro-koden . 
Någon ! Hallå ? 
Snälla ! 
Jag vet inte om nån ser det här , men om ni gör det ... 
Det var så dumt och jag är så ... 
Kyra , hör du mig ? 
Jag kommer in ! 
Hallå ? 
Jag är härborta ! Hjälp mig ! 
Mitt ben sitter fast . Jag vill inte dö ! Du kommer inte att dö . 
Jag lovar . Titta på mig . 
Jag drunknar inte . Jag har dig och ska få ut dig härifrån . 
- Tack . - Jag har dig . Allt är bra . 
Skåpbilen översvämmas snabbt . Vad händer ? 
- Är skåpbilens position säker ? 
- Jag vet inte . Den är upp och ner . 
Den åkte av vägen och hon sitter fast . Mår du bra ? 
Vad händer ? Prata med mig . 
Räddningsteamet kommer om tio minuter . 
- Det funkar inte . 
- Snälla , skynda er ! Kemi , vi måste ut härifrån . 
Jag tar fram bilder på hennes skåpbil . 
Det finns ett säkerhetslås på bakdörren till vänster . 
Kan du öppna dörren och dra ut henne ? 
- Jag kommer inte förbi sängramen . 
- Jason ? 
Hallå ? Hör ni mig ? Perfekt . 
Bara lugn . Kom här . 
Stanna hos mig . Jag lovar att få ut dig härifrån . 
- Snälla , jag vill inte dö . 
- Du kommer inte att dö . 
Vi gör det tillsammans . 
Du måste lita på mig . 
- Litar du på mig ? 
- Ja . Gör inte det , jag är galen . 
Allt kommer att bli bra . Det är bra . 
- Har du ett däckjärn ? - Nej . 
- Eller en kofot ? 
- Nej . - Har du ett rattlås ? 
- Det sitter nog under förarsätet . 
- Jag har det . 
- Hittade du det ? 
Bra . 
Det här kommer att funka . 
- Jag lyfter på tre . 
- Okej . 
Ett , två , tre . 
Herregud ! Tack ! 
Vi lyfter på tre . 
Ett , två ... 
Den rör sig ! 
- Mår du bra ? - Ja . 
- Varför tog det sån tid ? 
- Ingen orsak , sötnos . 
- Det här är kommissarie Batista . 
- Säg bara Nikki . 
- Jag vet inte hur jag ska tacka dig . 
- Kom här . Jag har sett så mycket av ditt liv att det känns som om jag känner dig . 
Det gör du på sätt och vis . 
Teddy gav aldrig upp hoppet en endaste sekund . 
- Det betyder mycket mer än följare . 
Kyra ! 
Jag trodde inte att jag skulle få se dig igen . 
Förlåt mig . Nej , förlåt mig . 
Jag borde inte ha blivit så arg . 
Om du vill att jag ska fria , så gör jag det här och nu . 
- Tack . För allt . 
- Givetvis . 
Njut av era resor . 
Jag hoppas att hennes möhippa är lite mer spännande än min . 
Vad menar du ? 
- Det blev inte vildare än så . 
- Du roar dig verkligen . 
Jag har haft galnare krogrundor . 
- Helen hade nog roligast av oss alla . 
- Jag ser det . 
Jag och Jay hamnade på en strippklubb . 
Japp . Vi blev uttråkade och drack några öl hos honom . 
Det var inte toppen alls . 
Förlåt om jag bröt mot reglerna . 
Händer det igen ersätter jag er båda med konstapel Hardbody . 
Han heter Jackson . 
Tror du att jag kan bjuda ut dig på en riktig dejt ? 
Jag vet inte . 
- Dejtar du alla dina klienter ? 
- Nej . 
Folk ser mig som ett sexpack till uthyrning och jag bryr mig inte om det . 
Jag faller för någons hjärna . 
Och du är så smart , Helen . 
Och bestämd . Du är min Elphaba . 
Fast jag skulle aldrig trotsa gravitationen . 
Det vore dumt , konstapeln ! 
Jag tror jag skadade handen . 
Jag vill bara lära känna dig . 
Om du låter mig . 
- Efter dig . 
- Okej . 
- Hej då . - Hej då . 
Åh , nej ! 
Tack , konstapeln ! 
Jösses ! 
" Jag är en dåre . Förlåt mig . 
Middag imorgon kväll ? " 
" Ett dussin rosor för varje timme mellan nu och då . " 
- Jag är redo för middag . 
- Ja , det är du . 
- Bara det inte är cheesesteaks . 
- Det blir det inte . - Bra . 
- Men vi kan dansa lite först . - Ja ? - Jag gillar det . 
- Gillar du det ? 
Jag gillar det inte , jag älskar det . 
- Är det inte Waynes ex ? - Har vi träffats ? Nej , men Wayne är min vän , och du måste fatta ett beslut . 
- Ursäkta mig ? 
- Jag har sagt min poäng . 
Okej . 
Städning . - Hej . - Hej . 
- Jag är lite upptagen nu . - Upptagen ? 
- Sträckkollar du Cartoon Network ? 
Jag är usel på att följa regler men ännu sämre med känslor . Känslor ? Jag bryr mig inte om känslor . 
Jag är bara trött på allt velande . 
Okej . 
Jag är ledsen att jag bara stack , jag kände mig bara så ... - Härinne ... 
- Som ett fångat djur ? 
- Ja , nåt sånt . 
- Jag tror jag fattar . 
Grejen är att jag tycker att vi är väldigt lika och jag antog att du skulle fatta varför jag är som jag är . 
- Jag tog med den här . 
- Han är redo för Gatorade . 
- Jag kanske inte är det . 
- Då är det min tur att vänta . 
- Men jag är väldigt törstig . 
- Jaså ? - Ja . - Hur törstig ? 
Väldigt törstig . Det är okej ... 
