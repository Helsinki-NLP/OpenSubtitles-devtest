" Tills lejonet berättat sin version , kommer jägaren alltid att vara hjälten . " 
När jag levde , var jag Cleo Johnson . Men som död , blev jag damen i sjön . 
Du sa att du visste vem som berövade mig livet , Maddie Morgenstern . 
IMORGON BEGRAVS " DAMEN I SJÖN " Du sa att ingen brydde sig innan du kom . 
Sanningen är att du kom i avslutningen av min historia och gjorde den till din inledning . 
Glad jävla postlåda . 
Okej . Tomtens lilla postlåda . Hepp ! 
Okej . Då så . Då kör vi . 
Hej , har du ett brev till tomten ? 
Glad thanksgiving , allihop . 
Med mig har jag Baltimores favorittv-värd , Wallace White . 
Vad tycker du om vår parad , Wallace ? 
Maryland Avenue är makalös , med gigantiska ballonger och allt . 
Titta på clownerna ! 
Wow . Och jonglören . Jag känner mig som en flicka igen ! 
Att vara barn på nytt är temat för dagen . 
Men oroa dig inte , pappa . Vi har nåt till dig också . 
Titta , här kommer våra Baltimore Orioles , som är ute på World Series-turné . 
Här kommer de dansande brevlådorna . 
Om ni nånsin har sett thanksgivingparaden , så vet ni att alla småttingar längtar efter samma sak . 
- Har du nåt brev till tomten ? 
- Och nu är stunden inne . 
Mannen som gör entré just nu kallas Sankt Nikolaus , tomten , den glade , men här i Baltimore kallas han jultomten . 
Stormande applåder när tomten äntligen anländer till Maryland Avenue , ända från Nordpolen . 
De tog med sig massor av gåvor och godsaker för de minsta . De kommer bli så glada . 
- Tessie . - Ursäkta . Tessie , kom . Här är pappa . Kom igen . Kom . Brexton är nog framkomlig . Har du nycklarna ? 
De är i din jackficka . 
- Hur vet tomten att vi är judar ? - Ja ? För att vi har en mezuza på dörren . 
- Och om jag sover över hos Mary ? 
- Han vet ändå . 
Mary skulle inte skvallra . 
Tomten finns inte på riktigt . Okej ? Marys feta pappa klär ut sig till tomte . 
Säg inte till Mary att din mamma sa så . 
Mary vet att han är fet . 
Pappa menar att säg inte till Mary att tomten inte finns . 
Jag är trött på att ljuga som en goy . Du är väl en stor flicka ? 
Om fyra veckor är det hanukka , då kan du be pappa om det du vill ha . 
- Okej ? - Jag vill ha en sjöhäst . 
Tills dess ... - ... får vi njuta av paraden . - En fin luch in kop . Här är också avstängt . Vi får gå tillbaka till Cathedral . 
Okej . Ge mig David . Kom . Du är en stor pojke . Varför parkerade du inte vid muséet som i fjol ? 
- Du sa att vi inte kunde parkera där ... - Nej ... 
En ögonätaralbino . 
Letar du efter nåt ? 
Jag bara tittade på fiskarna . 
Du borde komma tillbaka med dina föräldrar . 
Är de här ? 
Visste du att sjöhästar är fiskar ? 
Har du lärt dig det i skolan ? 
Jag går på Bais Yaakov . Vi lär oss inget om fiskar . Annat än att Gud skapade dem dag fem . 
Samma dag som fåglarna . Ja . 
Har du några sjöhästar ? 
Tebärstuggummi , tack . 
- Hej . 
- Mrs Schwartz . Bringa eller grytbitar ? 
Bringa för tre personer . 
Eller , för fem . 
Milton bjuder alltid in några i sista sekunden . 
- För att han är en sån mensch . 
- För att han är en macher . 
En macher vet vad som inte kan köpas för pengar . En vacker ayshes chail som springer och letar kosherlamm . 
Sex månader gammal . 
Oy , bara en bebis . 
Lugn , mrs Schwartz . Ingen kommer sakna honom . 
Ingen kommer sakna honom . 
Ursäkta . Får jag prova den gula klänningen i skyltfönstret ? 
Självklart , ma ' am . Ursäkta . 
Hon vill prova den gula klänningen i skyltfönstret . 
Självklart , ma ' am . Jag kommer strax . 
- Kan jag visa er nåt annat ? - Nej , tack . Det räcker med klänningen . 
Om hon inte hittar den i er storlek , kan jag beställa den . 
- Jag behöver nåt nu . - Då kommer den på måndag . 
- Jag lovar , vi hade tre i morse . - Och den i fönstret ? 
- Är ni säker ? Modellen är en ne ... - Det gör mig inget . 
Modellen har burit den hela morgonen . Den kanske är ofräsch . 
- Jag vill gärna prova den , tack . 
- Självklart , ma ' am . Jag följer er till provrummet . 
En dam vill prova den gula klänningen i skyltfönstret . 
- Gör det henne inget ? 
- Ethel för henne till provrummet nu . 
- Cleo . 
- Vi behöver klänningen . 
- Just nu , miss ? - Ja . Skynda . 
PROVRUM Stanna här . 
Klänningen har en svår hyska . 
Det är dragkedjan . 
- Hon kommer . 
- Jag får inte ner den . 
Jag kan göra det , miss Shirley . Får jag försöka ? 
Skynda . 
Är det därför gatan är avstängd ? 
En flicka från Pikesville är försvunnen . 
- Hennes föräldrar tog henne till paraden . - Åh , nej . Jag är från Pikesville . Jaså ? Det hade jag aldrig trott . 
Ni ser inte alls judisk ut . 
Hon dyker säkert upp snart . 
Det här är ju Baltimore , inte New York City . 
Tack så mycket . Jag tar kappan också . Tack . 
Nu sätter vi på dig nåt annat . Kanske en Mary Quant . 
Ursäkta . Klockan är redan tolv , och jag skulle få gå tidigt idag . 
- Det har inget sagt till mig . 
- Jag meddelade mr Goldberg förra veckan . 
Då får jag göra avdrag på din lön . 
Miss Shirley , kan jag få mina kläder ? 
Vänta . 
- Mrs Schwartz . 
- Tack , Aaron . 
Vad har hänt med din sko ? 
- Vad är det med din fåniga hatt ? 
- Allvarligt ? Jag ska ju hålla tal idag . 
Om hattar ? 
Du har bara den där hatten på dig så Myrtle får de rika vitingarna att tro att hon räddat lilla fattiga du . 
Eller så kanske hon anställer mig om jag ger ett bra tal . 
- Raring , du jobbar redan för henne . 
- Som volontär . RÖSTA FÖR KVINNLIGT LEDARSKAP 
- Ett annat ord för gratisarbete . 
- Du gör inte nog . Vår chef verkar ha bjudit in några av sina hejdukar . 
Säkert att du ska hålla tal åt Myrtle ? 
- Kan du inte vara snäll ? 
- Jag försöker . 
Den svart-judiska alliansen försvagas dagligen av Nation of Islams retorik om svart makt . 
Anti-semitismen är här för att stanna . Mamma . Trafiken . Hej . Hej . 
- Det var på tiden . - Förlåt . 
Är det här Seth ? Han växer snabbare än mina skulder . 
- Hej , mr Weinstein . - Maddie . 
- Milton , gör mig en toyve ... 
- Senare , Sid . 
Bara så du vet så är lägenheten i Sandtown tillgänglig igen . 
- Den i Bottom ? - Okej . En av dina killar fixade en hyresgäst i fjol . - Jag kommer till butiken ... - Det är thanksgiving . - Tack , raring . 
- Firar ni det ? 
- Det gör vi . 
- Inte jag . Vi är amerikaner . 
Förlåt att jag är sen . 
Allt är avstängd på grund av den försvunna vita flickan . 
Det här är min vän , miss Dora Carter . 
Givetvis , vi vet vem miss Carter är . 
- Ska ni sjunga för mrs Summer idag ? 
- Betalar hon ? 
Cleo , har du träffat Linda ? 
Hon är vicerektor på Douglas High School . 
- Vi möttes på charmskolans pristävling . 
- Jag donerade den där hatten . 
Jag hoppas få in min son Teddy i din skola . 
- Hans matteresultat är bäst ... 
- Hjälp mig välkomna Amerikas första svarta kvinnliga delstatssenator , ms Myrtle Summers . 
Och för våra priser , kallar vi upp vår vackra beskyddare , mrs Milton Schwartz . 
Tack , allihop . 
GE Jag vill tacka er alla och min make , Milton , för att du tillåter mig att representera vår familj idag . 
Vem behöver mig där framme när de kan titta på dig ? 
Jag vill tacka mina makalösa volontärer , de galanta damerna . Vissa av dem har varit med mig sen de bara nådde mig till knävecken , på den tiden jag undervisade . 
Som ni alla vet , tackar en judisk man Gud varje dag med de tre " She Lo Asani " - välsignelserna , för att inte ha gjort honom icke-judisk . 
Jag vet vad vårt samhälle behöver . 
För att inte ha blivit slav . 
En väg till välstånd . 
Och för att inte ha blivit kvinna . 
Man har sagt mig att det är på grund av de bördor vi kvinnor bär . 
Att skicka sina barn till fattiga skolor och bo i otrygga ... 
Våra skolor klarade sig bra tills er integrationslag skickade våra bästa elever till vita skolor . 
Han har rätt . 
Shell Gordon tycks ha skickat sina hejdukar för att störa eventet . 
Ingen har skickat mig . Jag talar för mig själv och affärsmän som mr Gordon , - som bryr sig mer om samhället ... - Affärsmän ? ... än ni gör . Mr Gordon är en brottsling som styrt det olagliga nummerlotteriet i 20 år , och nu lagt till droger till sin affärsmodell . 
Mr Gordon finansierade din första kampanj . 
Du för inte vår talan . 
Hon för min talan . 
Fortsätt , Cleo . 
Det här handlar inte om mr Gordon . 
Verkligen inte . Många av oss försöker bara se till att våra barn får en bra utbildning utan att behöva kämpa för att få en fjärdedel av det vita får . 
Som ni säger , vår värdighet kan inte tas ifrån oss . Den kan bara avstås . 
Jag är stolt att erbjuda detta pris till de tre kvinnor som personifierar syfte och ledarskap i vårt samhälle . 
Gratulerar , mina damer . 
Tack , mrs Schwartz . Jag har viktiga nyheter . 
Vi fick just veta att polisen lagt till en ny sökradie och en skallgångskedja kommer utgå var 45:e minut från Druid Hills synagoga . 
Delta gärna i sökandet och be för Tessie Durst och hennes familj . 
Lycka till . 
Jösses , mamma . 
Polisen har avsatt flera telefonlinjer . 
- Tessie Durst sågs senast ... - Jag borde ha åkt med pappa . - ... på en thanksgivingparad ... - Tessie Durst ? 
- Ja , Allan Dursts dotter . 
- Ja , jag vet vem Tessie Durst är . 
- Varför frågar du då ? - Jag frågar inte . Jag kan bara inte ... tro det . 
Jag kan inte laga mat . 
Vi borde leta efter henne . 
Mördade du Tessie Durst ? 
Det är lammet , Seth . 
Därför var jag sen . Jag fick köpa en ny klänning . 
Och du måste förresten laga mat , pappa bjöd in den där killen ni gick i skolan med , Wallace White . 
Det har han så klart inte berättat för mig . 
- Det var spontant . - Typiskt honom . 
Det var säkert spontant för Tessie Durst också . 
En liten judisk flicka försvann . 
- Vill du inte hjälpa till ? 
- Nej , jag vill äta . 
Om du försvann , skulle du då inte vilja att Allan hjälpte mig leta ? 
Så du vill leta efter Tessie så du kan räkna med familjen Durst om jag försvinner ? 
Varför är du alltid så arg på mig ? 
Lammet har legat i bilen hela dagen . Det är säkert skämt . Lammet är okej . 
Folk vill spela hos nån som hjälper dem välja nummer . 
- Vill du göra det måste du veta ... - Teddy ? 
Du ska allt få se . 
- Hur många gånger , Charlie ? 
- God eftermiddag , Cleopatra . 
- Charlie , du lovade mig . 
- Han delar Alvins talang för det . 
Shell höll inte på med droger när min pappa skötte lotteriet . 
Min son ska aldrig jobba för honom . Hör du mig ? 
Cleo , hur mås det ? 
Jag mår bra , Johnny . Kul att se dig . 
- Mamma , jag drar skämt . 
Jag vill ha mina kvinnor som solen . Strålande . 
Kul att se dig , Cleo . 
Du minns väl Eggy Woods och Johnny från Red Fox Lounge ? Japp . 
Glad thanksgiving på er . Kom igen , fortsätt du . 
Jag vill ha mina kvinnor som mitt kaffe . Hett och svart . 
Den där var bättre . Du börjar fatta grejen . 
Jag kan ett . Jag kan ett . 
- Hur går det där skämtet ? 
- Vilket ? Kom igen , Slap , du vet . 
Det där jag kommer hem och tror att ungarna är redo för thanksgiving . 
Gillade ni inte det skämtet ? 
Inte jag heller . 
Kom , gubben . Kom nu . 
Var så säker på att jag inte är klar med dig . 
Sluta , Leo . Eggy och Johnny kom just hit . - Dags att gå . - Det var åratal sen sist . 
Sätt på dig jackan , gubben . 
- Jag vet vad jag önskar mig till jul. 
- Du kan skriva ett brev till tomten . 
- Nej , han kan inte läsa . 
- Säger vem ? 
Teddy . Men jag ska rita en bild när min hand blir bra . 
- Varför sa du inte att hon var på väg ? - Har du ont i handen ? 
Sätt dig ner . Det är okej . 
Hans händer gjorde inte ont när han skrattade , - innan du kom in med din irritation . 
- Irritation ? Min irritation ? Du kan inte ens hålla Teddy borta från gatan . 
Teddy hänger inte på gatan . 
Grabben går ut varje dag och tar satsningar . 
Det skulle han inte behöva om ditt snuskiga nummer inte hade fått dig utkastad från varje klubb . 
Jag bor hos mamma tills du avgör om det är lika viktigt att börja jobba igen som att leva din sanning . 
Kom , Teddy . Vi går . 
Jag vet vem jag är och vem jag vill vara . 
Och hon är inte pank . 
- Det finns panka , lyckliga människor . 
- Är allt ett skämt för dig ? 
Pojkarna älskar mina skämt . 
- Knack , knack . 
- Vem där ? 
Hunden kissade . Hunden kissade vadå ? 
Hunden kissade på julgranen . 
- Såna skämt vill din mamma att jag drar . 
- Jag struntar i vilka skämt du drar . Bara folk betalar för dem , Slap . 
Kan du ta min handväska ? 
- Vänta , lämnar du mig på thanksgiving ? 
- Kom . 
Låt mig behålla en av pojkarna . Helst Teddy . 
Säg åt Shell att jag kommer förbi sen ! 
Du anar inte vad jag såg i bokaffären . 
På Highlandtown ? Ja . 
De två unga killarna som öppnat den , har startat en National States ' Rights Party-filial . 
De vill leka nazister . 
Leka nazister , alltså ? 
Det blir ingen lek om de startar en rörelse mitt i Baltimore . 
Stackars den jude som tror sig vara trygg . 
Jag tycker mer synd om lokala tv-stjärnor som inte har en dejt på thanksgiving . 
Tror du att kvinnor kastar sig över lokala nyhetsankare ? 
- Blygsamhet vinner du inget på . 
- Använd servett . 
Du kan väl presentera mig för några av dina vänner , Maddie ? 
- Tyvärr , Wallace . Maddie har inga vänner . 
- Det tror jag inte på . 
- Nej . Nån väntar alltid ... - Ska den ligga på golvet ? ... på att bli vän med Maddie Morgenstern . Förlåt . Schwartz . 
L ' chaim . 
Jag tog din mor till balen när Tessie Dursts pappa hade nobbat henne . 
Jag hittade henne tårdränkt i skolans nyhetsrum och tog ... Åh , Wally . Du är en sån historieberättare . 
Jag var inte tårdränkt . Jag grät . Och det handlade inte om nån fånig bal . 
Tänk om du hade gift dig med Durst . 
- Han har blivit alldeles för judisk . - Okej . Visa lite empati . 
Mannens dotter är försvunnen . Knappast läge att skämta om honom . 
Jag har aldrig hört talas om denna skolflickskärlek till Allan Durst . 
För att det var ingen skolflickskärlek . 
Jag var upptagen av skoltidningen mitt sista år . Det var allt jag brydde mig om . Ingen såg mig ens . 
Vem är blygsam nu ? 
Alla var förälskade i henne . 
Men bara Milton hade den hemliga ingrediensen . 
Det räcker . Säg inte sånt framför Seth . 
Ska skoltidningens stjärna äntligen kolla till lammbringan ? 
Bra där . 
- Ja , mycket bra . - Han har tv-utseende . 
Visst har han ? Det säger jag till honom . 
När vi kommer hem lägger vi kalla kompresser på dina händer . 
Det dämpar svullnaden . Då kommer du må bättre . 
Förlåt . Förlåt mig . Lägg in den där påsen åt mig . 
Jag vet , raring . Jag vet . Ja . 
Jag vet . Låt mig ta av den här . 
Jag vet . Hej , mamma . 
- Här . Kom och sitt med mig . 
- Var är Slappy ? 
Han ska jobba . 
Då måste du ha hittat en ny man . 
Glad thanksgiving . 
Den vore gladare om du tillbringade den med familjen istället för bakom baren . 
När mrs Summer ger mig heltid slipper jag jobba kvällar . 
Jag behöver bara lite hjälp med pojkarna tills dess . 
Bara över helgerna . 
Bara om ni alla klämmer in er i ett rum . 
Hur mår min lilla gubbe ? Kom . Låt mig få titta på dig . 
- Hans ögon är gula igen , Eunetta . - Jag vet . - Han har läkartid imorgon . Lite juice ? 
- Han har fått nog av läkare . De säger bara att sicklecellsjukdom är obotlig . 
- Mamma ... - Profeten måste komma och kika på honom . 
- Skit i profeten . - Hallå . 
Tänk på språket . 
- Du hörde . Han rör inte min son . 
- Tänk på vad du säger om pastorn . Tänk själv , Isaiah . 
- Du verkar glömma vems hus du är i . - Vadå , min fars hus ? Den stafettpinnen tog jag över för länge sen . 
Du sitter bra i hans stol . 
Du ska visa Isaiah respekt när du pratar med honom . 
- Respekt går åt båda hållen , mamma . - Det tål att upprepas . 
Jag måste till jobbet . 
Lägg lite varma kompresser på hans händer och ... 
Kapten Stassley hos Baltimorepolisen har meddelat att han gett flera enheter i uppgift att söka efter flickan , och har sagt åt alla patrullerande poliser att hålla utkik efter misstänkta . 
Tessies försvinnande har enat en stad som alltför ofta varit kluven . 
Biskop Carol och pastor ... Allan Durst . 
Vem bryr sig ? 
Om ni har information som kan hjälpa situationen ... Är det nåt mer du vill säga ? 
Tessie Durst är försvunnen . 
- Det känns fel att stå i köket just nu . 
- Jag trodde du gillade det nya köket . 
Maddie , kan vi inte bara njuta en trevlig thanksgivingmiddag utan att prata om Tessie Durst i några timmar 
Mr Durst , vill du säga några ord till våra lyssnare ? 
Snälla , be för vår älskling , och håll utkik efter henne . 
Vi håller hoppet uppe och väntar på att få hem henne igen . 
- Maddie ... 
- Vi borde göra dem sällskap . 
... du använde mejerifaten till bringan . 
Varför gjorde du så ? 
Jag beklagar , allihop , men jag måste kasta bringan . 
- Förlåt , Wallace . - Ingen fara . - Förlåt Wally ? - Förlåt ... Ja . Åkte Wally ända till Lombard Street för att köpa kosherlamm ? 
Wallace är vår gäst , och nu har vi inget att servera . Eller ska vi vänta tills de hittat Tessie Durst innan vi äter ? 
Visst . Vi kan fasta . 
Jag trodde det var thanksgiving , men det är väl Yom Kippur . 
Vad gör ... Hallå ... Ge mig den där . Vad gör du ? 
Ge den till mig . 
Ursäkta mig . 
Vad ... Wallace har gått . 
Kan du komma ut och sluta med galenskapen ? 
Jag har städat undan allt . 
Kom , låt mig få se på din hand . 
Vad är det ? Vad har det tagit åt dig ? 
Varför beter sig alla som om det är fel på mig för att jag bryr mig ? 
Om Tessie Durst ? 
Jag vet inte , Maddie . 
Hela Baltimore letar efter henne , men jag är en meshuggener ? 
Jag vet ingen annan som reagerar på det här sättet . Och jag sa aldrig meshuggener . 
Det sa jag inte . 
Jag var bara upprörd över att vi inte hade nåt att servera . 
Okej ? Gud förbjude att det går en dag utan att jag betjänar dig . 
- Betjänar mig ? 
- Ja , Milton . 
Ja , Milton . Jag har tjänat dig i 20 år . 
Och du tycker inte att jag duger till nåt annat än hemmafru . 
Det gör jag inte alls . 
- Jo . 
- Nej , det gör jag inte . Nej . 
Vad är det då ? Maddie ... Vad tycker du att jag duger till ? 
Du har aldrig velat göra nåt annat . 
Jag försökte aldrig göra nåt annat ! 
Har du aldrig undrat varför ? 
Om ett saknat barn inte hittas inom de första 24 till 48 timmarna , är barnet förmodligen dött . Har du hört det ? Maddie , vad är det här ? Vad är det här ? 
Vad är det som pågår ? 
- Låt henne gå för fan . - Tänk på språket . 
Jag behöver inte din fars tillåtelse att gå . 
Svara mig , Maddie . Vart är du på väg ? 
Vad är det som pågår ? 
Maddie , det här kommer från ingenstans ! Helt från ingenstans ! 
En gång i tiden hade jag inte trott att du skulle lämna din man , ditt fina hem , livet ni hade tillsammans . 
Men precis som döden förändrade hur folk såg på mig , förändrade det hur jag ser på dig . 
Jag såg dig , Maddie Schwartz . 
Innan allt det här började , så såg jag dig . 
Jag såg dig se mig se dig . 
Det är som en tungvrickare man säger som barn . Jag målade en tavla av mig som målade en tavla av mig som målade en tavla av mig . 
Och så fortsätter det tills allt blir så smått att man inte ser nåt alls . 
- Godkväll , mrs Johnson . 
- Hur mår Dora ? 
Svartpeppar och varmt vatten kanske hjälper . 
Jag tittar till henne när jag är klar . 
- Hänger du in den här ? - Självklart . Tack , Clarence . 
Den försvunna flickan fick judarna att stänga tidigt . 
Du vill att jag säger till mr Gordon att vi inte har nån försäkring när hela staden satsar på 466 ? 
Leo , glad thanksgiving . 
- Glad thanksgiving , Vernon . - Ja . 
Jag kommer . 
- Vad gör du här ? Kom in . - Sid , förlåt att jag stör . Kom . Det är inget besvär . 
Lägenheten du nämnde , den i Bottom . - Jag vill befria dig från den ett tag . 
- Vad pratar du om ? 
Var är Milton ? Vi har stängt . 
- Men vi har ... 
- Kom hit med den . 
Tack , grabbar . 
Stackars Tessie . 
- Dra åt helvete . 
- Det är Cleo . 
Förlåt . 
- Dra åt helvete , Cleo . 
- Du uppträder kl 22 : 00 ikväll . 
- 23 : 00 . 
- 22 : 00 . 
Jag tog med pepparvatten . 
Har du fortfarande den dumma hatten på dig ? 
Fan ta dig , Dora . 
Vad har hänt med din hand ? 
- Ska jag sluta ställa frågor ? - Det skulle uppskattas . 
Jag kan be Judith visa dig lägenheten . 
- Minns du min dotter ? Judith . - Självklart . 
Judith ! Ja ? 
Jag vill att du visar lägenheten för mrs Schwartz . 
- Den i Bottom ? 
- Hur många lägenheter har vi ? 
Skärp till dig . 
Maddie , det är ingen brådska . 
Jag köper tillbaka dem . Jag ska bara panta dem en månad eller två . 
- Den är inte köpt här . 
- Han köpte den på Steiner ' s. 
Steiner ' s. 
Snobbigt värre , men nu har de stängt . 
Vad är det jag brukar säga ? 
" Man behöver inte kristallkronor för att sälja diamanter . " 
Just det . 
Jag kan bara betala 500 . 
Men Milton har försäkrat den för 2 000 dollar . 
Så här gör vi . Jag vill inte hamna i kläm här , men om nån kommer in och vill ha den här stilen , så kan vi komma överens . 
- Hittade du nycklarna ? 
- Jag kollar där bak . 
Här . 
Jag väntar i bilen . 
Och Maddie ... Glad thanksgiving . 
- Vad händer , Curtis ? 
- Bara en vanlig kväll på Pharaoh . 
- Är det full fart ? - Ja . 
Hur går det här ute ? 
Inte alls . Jag borde nog komma in . 
Jösses . 
Det är bara för klubbmedlemmar . Det vet du . Du borde testa kuddkrig . 
Bara klubbmedlemmar , sa jag . Det vet du . - Och artister . 
- Du uppträder inte här längre . 
Har Shell sagt det ? 
Pratar du med mig pratar du med mr Gordon . 
Mannen , jag bad Cleo säga till Shell att hennes make skulle komma förbi , okej ? 
Jaså , det gjorde du ? 
Vänta här ute om du vill . 
- Har nån av er sett Shell ? 
- Mr Gordon är på scenen . 
Ge en applåd för mannen , munnen , myten , Roy " Tanglefoot " McCoy . 
Chefen , Slappy är där ute . Han vill göra ett set eller nåt . 
- Vill han ? - Ja . Jag vet inte vad jag ska säga . Säg åt Cleo . Visst . Okej , chefen . 
Konstapel Platt . 
Reggie , hur är läget ? 
Ditt på det torra ? Inga dumheter ? 
Hela dagen , varje dag . 
Nån har gett dig en blåtira . 
Jag tar dem nästa gång . 
Slappy vill komma in . 
Vad glor konstapeln på ? Borde inte du leta efter den försvunna flickan ? Innan de kommer hit och spöar våra bröder ? 
Mitt skift börjar om en timme . 
Ska jag hitta henne , måste hon fortsätta vara försvunnen till kl 22 : 00 . 
Eller hur , Reggie ? 
Snabb service innebär inte att du slipper ge dricks . 
- Jag ger dricks . 
- Inte tillräckligt . 
Jag visste inte att min lilla paus skulle orsaka sånt besvär . 
Jag skulle inte kalla det paus när du inte är i tjänst . 
Ers nåd , försöker jag visa mig oskyldig till att vara snål eller menar du att jag tar mutor ? Jag undrar bara vad du gör här mitt i veckan . 
Samma som alla andra . Musiken och utsikten . 
- Utsikten ? - Ja . 
Oroa dig inte för mig . Jag kissar inte på tjingade träd . 
- Jag visste inte att du gillade träd . 
- Varför skulle jag inte ? 
Svårt att hitta vita träd . 
Dora . Dora ! 
Blomster med konster ! 
Dagsslutsrabatt ! 
Köp medan ni kan . 
Revolutionära jordgubbar färskare än Martin Luther King . 
Blomster med konster ! 
Köp medan ni kan ! 
Dagsslutsrabatt . 
- Låt mig hjälpa dig . 
- Tack . 
Ja . Det här är så trevligt . Ska jag skaffa en hopvikbar säng ? 
Det enda sättet mamma släpper ut mig ur huset utan en man är om jag flyttar in hos en trevlig kvinna från Northwest Baltimore . 
En trevlig äldre dam . 
Jag har inte ens sagt till min mamma att jag lämnat . 
Det kommer inte bli lättare än när jag var 20 . 
Så gammal är du inte . Och får jag flytta in hos dig slipper du panta din ring . 
Är vi nära ? Ja . Det är hitåt . 
Kom . 
Vad gör du där borta , pinglan ? 
Dörren bara fastnar . 
Den där fungerar inte . 
Det här är badrummet . 
Badkaret är rätt stort , vilket är trevligt . 
Det är lite lortigt för jag råkade lämna fönstret öppet . 
Han blev sur på mig för det . 
Ja , men ingen har bott här på fem , sex månader . 
Jag hade tänkt att jag kanske skulle flytta in , men det var mitt fel . 
Jag kan komma tillbaka med en svamp eller en mopp om du vill . Och en kudde . 
Ja , jag verkligen ... Jag älskar den här lägenheten . Jag har alltid velat bo här , men pappa vägrade . 
Han blir så orolig för mig . 
Jag vet inte vad du tycker om att dela , men jag har inget emot att sova på golvet . 
Jag tar den . 
Jag ska hjälpa dig med din väska . Nej . Tack . Jag ska bara byta om , sen går jag till synagogan och hjälper till med skallgångskedjan . De låter inte en kvinna vara med . 
Då startar jag en egen kedja . 
Det är ingen kedja om du går ensam . 
Jag vill inte ha en rumskamrat . 
En vän då ? 
Vad är det ? 
- Kom igen . Upp . - Nej . Dora . Dora . Jag svär , om du inte är på scenen om tio minuter ... Kom igen nu . 
Så ja . Kom igen , baby . Din chef fick henne att börja . Hur ska hon kunna sjunga ? 
Min chef ? 
Är inte du här ? - Du jobbar också för honom . 
- Jag gör inte sånt du gör . 
Kom igen , baby . Cab Calloway kommer ju ikväll . 
Så ja . 
Din jävel . Här . Du vet ju att mr Hi-De-Ho vill höra dig sjunga . 
Ta ut henne på scenen när hon öppnat det andra ögat . Det dröjer inte länge . 
Så ja , baby . Mr Hi-De-Ho längtar efter att höra dig sjunga . 
Lefty , Dora går på om fem . " Where Did Our Love Go , " halvtempo . 
Cleo . 
Shell . 
Ville ni prata med mig , mr Gordon ? 
Ja , sätt dig ner . 
Vill du ha en drink ? 
Nej , tack . 
Cleo har skött mina räkenskaper sen hon gick i ankelstrumpor . 
Dessutom jävligt bra . Jag försöker ge henne mer jobb , men hon är för upptagen av att hålla tal . 
Eller hur , Cleo ? 
Du är kallsinnig . Lämnar Slappy där ute som en gammal hatt . 
Ja , vi har haft en tuff dag , och jag ville inte ta med den hit . 
Jag vill inte se ännu en svart man misslyckas , så vi låter honom göra ett set . 
- Tack , mr Gordon . 
- Jobbar du med mrs Summer nu ? 
Nej , jag jobbar som volontär 
- för mrs Summer . - Så du jobbar gratis ? Och jag betalar för ditt arbete ? 
- Nåt gör jag allt fel . 
- Det gör du . 
Du kan väl gå ut på scenen och berätta för snubbarna att Dora kommer förbluffa dem . 
Jag ogillar strålkastarljus , mr Gordon . 
Kom ihåg det nästa gång mrs Summer ber dig hålla tal . Det är skillnaden mellan henne och mig . 
Jag betalar dig , så det är en order . 
Ja , sir . Ursäkta mig . 
Duktig kicka . 
Tessie ! Tessie . 
Jag vet vart jag ska . 
Det finns en stig här nere som leder till sjön . 
Är det här ditt gamla hångelställe ? 
Nej . 
- Varför beter du dig så skumt ? 
- Det gör jag inte . Okej . 
Det är faktiskt inget fel med att rulla naken i gräset med ett par pojkar . 
Kan du hålla den här ? 
Det är 1966 . 
Jag rullade inte naken i gräset med nån . 
Vad gör du ? 
- Vad ser det ut som ? - Rök inte nära mig . 
Mina damer och herrar . Nästa sångfågel har jag känt sen jag var en liten flicka , och jag vet ändå inte vad hon ska göra härnäst , men hon får mig alltid att vilja ha mer . 
För ert höga nöje , den unika och oförglömliga miss Dora Carter . 
Det är fan inte sant . 
Vänta ! 
Rör henne inte ! 
Jag vill hålla om henne . 
- Bara ... - Håll om mig . 
Judith , gå och hämta hit nån . 
Jag lovar att inte röra henne , men jag måste vänta här med henne . 
Om du vore mor skulle du förstå . 
När man dör , är man inte en flicka längre . Eller en kvinna . Eller en maka . 
Man är ingens moder , ingens dotter . 
Och ingen kan säga åt en hur man ska leva sitt liv . 
Du ville väl att Tessies död skulle göra dig fri ? 
Men den visade dig bara till dörren . 
Min död fick dig att öppna den . 
