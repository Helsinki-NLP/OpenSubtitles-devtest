Ruby ! 
Ruby ! 
Din väckarklocka har ringt i tio minuter nu . 
Förlåt att jag väckte dig . 
Du såg ut att drömma nåt trevligt . 
Fin hoodie . 
Göm den för mamma . Om hon tvättar den försvinner lukten . 
Närhet och avstånd utesluter inte alltid varandra . 
Man kan känna sig nära människor som är långt borta , eller lita på nån som man ogillade för bara två veckor sen . 
Tack för igår . 
Det var verkligen snällt av dig och ... 
Tack för igår . Du behövde inte köra mig ända hem . 
Jag trodde mig veta hur man tappar kontrollen . 
Alkohol , sex , droger . 
Jag insåg inte att det bara är lekar . 
Igår fick jag uppleva att tappa kontrollen över mina känslor . 
Tack . 
- R.J.B. 
Du har aldrig berättat vad J står för . 
Och det kommer jag aldrig göra . 
JAMES Erkänn att det står för James . - J.M.B. 
Självförtroendet i topp , verkar det som . 
Du undviker frågan . 
Måste vara nåt hemskt . 
Jag berättar om du avslöjar ditt M ? 
Snyggt försök . - J.M.B. 
Mår du bättre nu ? 
Ja ... Men jag är nervös för idag . 
Oroa dig inte . 
De flesta såg bara min blöta rygg igår kväll . 
Då hade de i alla fall en trevlig kväll . 
Ruby Bell , försöker du flirta med mig ? 
Maxton Hall THE WORLD BETWEEN US 
EFTER ROMANEN " SAVE ME " AV MONA KASTEN 
Bagarens dotter ... 
Varför stirrar du ? 
Alla tittar på mig . 
Bry dig inte om det . 
Tillämpa Beaufort-koden : Total nonchalans , oavsett situation . 
Du ser ut att behöva en örfil . 
Jag kanske gillar örfilar . 
Är det där Ruby Bell ? 
Hon är cool och nonchalant . 
James Beaufort bar henne i sina armar . Vilken lyckost ! 
- Sluta ! Eller , äsch . - Utmärkt . 
Efter lite övning tror du på det själv . 
Tro mig . - Maxton ! - Hall ! 
Du saknar det , va ? 
Kom igen , män ! Vi är vinnare . 
- Vi är vinnare ! - Till skillnad från dem . 
ELAINE Ring mig ! 
Lydia , sluta ignorera mig och svara . 
Är han ihop med socialfallet ? 
God morgon . 
Vill du ha en kanelbulle ? 
De kommer från bageriet i Compton . 
Tack . 
Jag måste tacka dig . 
Utan dig skulle vi inte ha en ny kollektion imorgon . 
Det finns så mycket passion och kreativitet i hela konceptet . 
Innovation . Kvalitet . 
Allt som Beaufort representerar . 
Och allt det måste James förkroppsliga imorgon . 
Vad vet du om den här tjejen ? 
Ingenting . 
Hon går visst i vår skola . 
Det var bara ett dumt festskämt . 
Några skojade i poolen . 
Att bli involverad med fel person kan förstöra ens liv , det vet ju du . 
Jag fick betala ditt ex 500 000 pund för att förstöra fotona han hade . 
I morgon ska din bror bana väg för er båda . 
Young Beaufort är bara början . 
Nästa kollektion kanske bär ditt namn . 
Du kan klara det . 
Men nu är det viktiga att James inte förstör presskonferensen . 
Han får inte tappa fokus . Inte nu . 
Ni står nära varann . 
Använd det . 
James . Vet du vem jag åt frukost med i morse ? 
Pappa . 
Du måste vara försiktig med Ruby . 
- Bad han dig att prata med mig ? 
- Ja , typ . 
- Det är bara ett foto . - Bara ett foto ? 
Om han tror att du är distraherad blir det ett himla liv . 
Jag har koll . 
- James . - Lydia . 
Det är bäst att du skärper dig . 
- Annars ingriper han . - Oroa dig inte . 
Ruby är åtminstone ingen lärare . 
- Lådorna är för tunga för dig . - Kan vi hjälpa dig ? 
Nå , hur var han ? 
Är det sant vad de säger ? 
- Vadå ? 
- Du vet . 
Gjorde ni det ute eller i hans limousine ? 
Säg att ni gjorde det i limousinen . 
Det lämnar jag åt er fantasi . 
Och ljusen ... 
- Alla tror att jag har legat med James . - Och ? 
Nej . Vi har inte ens kysst varann . 
Han räddar ditt liv , dumpar sina vänner , och bär iväg med dig som Miss Wet T-shirt , i månskenet , men kysser dig inte ? 
Vad mer behöver ni ? Fyrverkerier ? 
Videorna är uppladdade överallt . 
Om du dejtar en kändis , får det uppmärksamhet . 
- Men var det en dejt ? - Ville du det ? 
Hej , Ruby . 
Den frysta maten levereras snart . 
- Isbitar , kött ... - Tack , Kieran . 
Lugn , jag tar hand om det . 
Ta hand om bordet också . 
De ska vara därinne . 
Vad har du gjort med den stackaren ? 
Han gör sig inte till för mig . 
Fast det är sexigt . 
En man kan vara artig mot en kvinna utan baktankar . 
Jag är inte helt säker på att Rutherford är en man . 
Tack . 
Den första skolfest jag sett fram emot . 
Kanske jag t.o.m. kommer i tid . 
Då hinner du till Rubys födelsedag . 
Är det imorgon ? 
Visste du inte det ? 
Lexington ordnar ett kalas åt mig . 
Då kommer jag definitivt i tid . 
Vem ska du annars dansa första dansen med ? 
Det finns säkert nån . 
Ruby ... Du ville att maten ... Den skulle vara så färsk som möjligt , eller hur ? 
Vi kan slakta dem själva . 
Ska vi slakta 150 rapphöns i skolköket ? 
Självklart inte . 
Ruby , jag fixar det . 
Jag kanske kan ... 
Burarna måste bort . Nånstans där det finns frisk luft . 
Ni hörde Ruby . 
Bra . Mr Lexington , jag har en fråga om ... 
Och Rutherford . 
Bra jobbat . 
" Bra jobbat . " 
- Som hon ser på honom ... 
- Ja , de har varit ihop ett tag . 
Har de ? 
Ligger du med henne ? 
Vad ? 
Eller återupplivar ni bara gamla minnen ? 
Ni jobbar tillsammans . 
Det kan vara extremt praktiskt eller extremt besvärligt . 
Vill ni fråga om provet vet ni var jag finns , miss Beaufort . Men nu måste jag gå . 
Är det så lätt för dig ? 
Att återgå till det gamla ? 
Att bara vara min lärare igen ? 
Var det inte planen ? 
Att låtsas som om inget hänt ? 
Du ser ju hur glad ut som helst . 
Hur ska jag se ut ? Som om jag förlorat min stora kärlek ? 
Se inte på mig så där . 
Varför inte ? 
Då kanske jag gör nåt jag svurit på att inte göra igen . 
Lydia . Vi måste hålla oss till planen . 
Strunt i planen . 
Vi ger oss av . I dag . 
Vi börjar om nån annanstans . 
Byt jobb . Jag tar examen . 
Det vill du inte . Inte på riktigt . 
Lämna ditt hem , din familj , dina vänner . 
- Jag vill vara med dig . - Inte så . 
Jag gör inte så mot dig . 
Du vet inte vad jag vill . 
Men du är tydlig med vad du vill . 
Hur mår Ruby ? 
Bättre . 
Bra . 
Cyril är en stor idiot . 
Det är inget nytt . 
Det var en händelserik kväll . 
Ursäkta att jag klampade in . 
Kesh såg inte jätteglad ut . 
Nä . 
Han är inte redo . 
Hur funkar det för dig ? 
Jag är jättekär . 
Det hjälper . 
Tänka sig att få se James Beaufort dra 600 vaktlar över gården för ... En tjej ? 
Det är rapphöns , inte vaktlar . 
Och du får gärna hjälpa till . 
Visst . Vart då ? 
Nånstans i friska luften . 
" Och därför är det min stora ära ... 
" Mitt stora nöje och en ännu större ära , " att följa i mina föräldrars fotspår " och presentera den nya kollektionen som junior-vd . " 
- Öva på det . - Ja . 
Hur var coachningen med Charles ? 
Har du några frågor ? 
Självklart . 
Du är förstås väl förberedd för den viktigaste händelsen i ditt liv . 
Du har studerat mina mejl i flera dagar , antecknat alla datum noga , lärt dig alla ord utantill , och studerat den nya kollektionen i minsta detalj . 
Jag vet vad som väntas av mig . 
Imorgon , James , blir du mr Beaufort ... Junior . 
Jag har bjudit in PR-chefen på middag efter presskonferensen . 
Var redo . 
Men jag måste till galan för donatorerna . 
Livet handlar om beslut , James . 
Och vet du varför ? 
För att vi inte kan få allt . 
Förälskelse gör oss till idioter . 
Vad väljer du ? 
En förälskelse du har glömt om två år , eller din familj ? 
Det är ditt beslut . 
Men det är jättebra om du kommer . 
Så att vi kan fokusera på det viktiga . 
Har den äran idag 
Har den äran , kära Ruby 
Har den äran idag 
Önska nåt ! 
Nå ? Är det rätt ? 
Nämen , Gud ! Tack , pappa ! 
Del fyra i Förberedelser för Oxford . Nu fattas bara del fem . 
En tegelsten till . Hurra . Öppna min nu . 
Nämen ! Del fem . Vilken överraskning ! 
Tack . 
Får jag äta tårta nu ? 
Sakta i backarna . 
Här är en present till . 
- Visa . Vad är det ? - Den är min . 
- Visa mig . - Nej . 
Måste till skolan ! 
Vem går i skolan en lördag ? 
- Mamma , hjälp mig . - Ja . 
Nej , vänta ! 
Förlåt för det jag sa . 
Du hade rätt . 
Jag ville bara tro att det är jag som bestämmer över mitt liv . Inte han . 
Det är orättvist . 
Vad vet du om orättvisor ? 
Pappa pratar bara med mig för att utpressa mig . Mannen jag älskar ligger med sitt ex och du får presentera konceptet som jag jobbat med i åratal . 
Allt jag bryr mig om är antingen inte mitt , eller fel . 
Du vet inte hur det är att vara allas reservplan . 
Gör oss båda en tjänst och spela din roll . Det blir bäst så . 
Vi kanske kan byta , som i Föräldrafällan . 
Du tar presskonferensen , jag galan . 
Jag kan ha lösmustasch . 
- Ingen märker nåt . - Aldrig . 
Allt bra ? 
Pappa har bjudit vår PR-ansvariga på middag . 
Jag missar galan i Maxton Hall . 
Och Rubys födelsedag . 
Evenemanget är viktigt för företaget . För pappa , mamma och Lydia . 
Det känns skitjobbigt . 
Det är bra . 
Smärta är en signal att du är redo för förändring . 
De är överallt . 
De andra fångar dem . Dekoratörerna kommer snart . 
Hur ska de kunna jobba med tusen fåglar runt sig ? 
- Bara 150 . - Upptäcker Lexington det , är jag körd . 
Körd . 
Då så , vad väntar du på ? 
Och grattis . 
- Här bakom . - Okej . 
Låt den inte smita ! Fan ! 
- Säkert att den är härinne ? 
- Ja . De är väldigt snabba för att ha så små fötter . 
Som du . Det kanske var så du fick ditt mellannamn . 
Jag tog reda på det som jag lovade . 
Jemima betyder " duva " . Det är ett gulligt namn . 
- Ser du den nånstans ? 
- Nej . 
Paus ? 
Paus . 
Tack för presenterna . 
Väskan är jättefin . Och teckningen ... 
Tänker du avslöja ditt mellannamn nån gång ? 
Jag kan brodera det på nåt . 
Jag har fullt upp med märkta kläder , tack . 
M står för Mortimer . Efter pappa . 
Jag kommer inte ikväll . 
Vi lanserar vår nya kollektion och pappa vill att jag träffar PR-personen . 
Jag är ledsen . 
Det blir säkert kul . 
Jag vill bara få det överstökat . 
Jag vill inte gå på presskonferensen eller ta över Beaufort . 
Jag vill kanske inte ens gå på Oxford . 
Menar du det ? 
Du hade rätt på förberedelsekursen . 
Jag är inget mer än mitt namn . 
I teorin har jag en massa privilegier och möjligheter , men ... Inget av det är mitt beslut . 
Och vad vill du ? 
Vad skulle göra dig glad om du fick göra vad du ville ? 
Jag vet inte . 
Jag tror att alla har stunder när de glömmer allt omkring sig . När de slutar ifrågasätta varje steg och tanke och bara följer sin instinkt . 
Livet handlar om att tillåta den tanken . 
Och ta reda på vad man brinner för . 
Jag fick tag på den sista . 
Bara så att jag förstår , miss Bell . 
Först säger ni att han förstörde er fest , sen vägrar ni arbeta med honom , nu ber ni mig att korta av hans straff - och låta honom spela lacrosse igen ? 
- James hjälpte till med festen , han hittade på temat och genomförde det . 
Han har förstås gjort dumma saker förut , men nuet är det som betyder nåt . 
Om denna fest blir lyckad , som den blir , är det tack vare honom . 
- Okej . - På riktigt ? 
Ja . 
Om festen avlöper utan problem , - får han spela igen . - Tack , sir . 
Men , miss Bell ? Glöm inte vad mer som står på spel ikväll . 
Inte bara för mr Beaufort , för er också . 
Pappa ska ta hem rapphönsen till vår gård . 
Vi ska få hit kyckling istället . Som inte lever . 
- Ursäktar du mig ett tag , Kieran ? - Ja . 
Stor kväll . DONATIONSGALA 
Inte bara för mig . 
Ska jag skicka några strippor ? 
Gå din väg . 
Se till att få din rekommendation . 
" Idag börjar ett nytt kapitel för oss alla . " Därför är det ett stort nöje och ... " 
" En ännu större ära att följa i mina föräldrars fotspår " och presentera vår nya kollektion som junior-VD . " 
Otroligt att du kan talet utantill . 
Jag skrev det ju . 
" Men oroa dig inte , James banar väg för er båda idag . 
" Nästa kollektion kanske bär ditt namn . " 
" Livet handlar om beslut , för vi kan inte få allt . 
" Vi behöver dig . " 
Det slutar aldrig . 
Det finns alltid nåt viktigare än vad vi vill . 
Tills det är vi som bestämmer . 
Få motståndaren att tro att den bara har en möjlig utväg . 
Percy . 
Vänd om . 
Låt dem inte stöta på dig eller tafsa . 
Ta en taxi hem , vi kan inte hämta dig . 
Jag ska . 
Jag har en idé för ditt hår . 
Raring ? Ha så kul nu . 
Tack . 
Ruby , kan du inte chilla i fem sekunder ? 
Jag chillar . 
Vi har slitit hårt med den här festen . 
Och se dig omkring . Det är perfekt . 
Du fyller år idag , och är jättesnygg . 
Du får din rekommendation , vi åker till Oxford och blir politikens Beyoncés . 
Och du är en prinsessa även utan din prins . 
Så kan vi njuta av kvällen nu ? 
Vad har vi blivit ? 
Smartphone-zombier . 
Sluta kolla din mejl . Fixa dejter . 
Här är en . En till . Vad heter appen ? 
Nu ska vi hitta din drömprins . 
Titta , vad söt . 
Han då ? 
Snyggare än jag . 
Skulle du nobba mig också ? 
Du är bara sur för att Lydia bangade . 
Det gjorde hon inte . 
Hon dök bara inte upp . 
- Exakt . - Jag vet inte . 
Om Alistair inte finner lyckan , måste vi hjälpa honom . 
Vi hittar nån till honom . Vad sägs om honom ? 
Eller honom ? 
Sluta . 
Sluta med den här toxiska maskuliniteten . 
Säg bara vilka du tycker är snygga . 
Sluta nu ! 
Den här är bra , fast ansiktet syns inte . 
Är det ett problem ? 
Föredrar Alistair knubbiga män eller mer maskulina och muskulösa ? 
Vad vet jag ? 
Jag är helt straight . 
Jag har en match . 
Man kan tveka hela livet . Men bara om man hoppar får man veta vad som finns utanför klippan . 
En avgrund ? Eller en bärande vind ? 
Att förlora fotfästet är skrämmande . 
Om man fokuserar på sina drömmar glömmer man att tyngdkraften kan lura en . 
Ibland är det handlingen . 
Att man genom att ta sitt öde i sina egna händer kan bli nån annan . 
Var fan är James ? 
Där han ska vara . 
Precis som jag . 
Vad gör du här ? 
Vi har tre timmar kvar av din födelsedag . 
Vi borde njuta av dem . 
Jag har en överraskning åt dig . 
Jag pratade med Lexington . 
Om festen går som han vill får du spela lacrosse igen . 
Vad ? 
Ruby Jemima Bell . 
Måste vara en säkring . 
Proppskåpet är i västra flygeln . 
Det var ditt sista uppdrag i kommittén . 
Det var kul att jobba med dig . 
Det låter som att du säger adjö . 
Är det så här det ser ut när du vet vad som förväntas av dig ? 
