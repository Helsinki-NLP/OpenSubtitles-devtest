- Åh , herregud , vad ? 
- Jag kollade precis ditt schema . Du tycks inte vara upptagen just nu . 
Jag är nervös inför provspelningen . Vill du öva repliker med mig ? 
Okej . 
Dustin vill ... skapa förändring . 
- Göra skillnad . - Javisst . Amerika är ganska rörigt . Det är orättvist att det inte finns nog med paj så att alla får sin bit vid bordet . 
Och du har arrangerat en hel presskonferens för att meddela detta . 
En enorm presskonferens . 
Nåväl , jag ser fram emot det . 
- Julio , hon är här . - Förlåt , jag måste gå . 
Jag har en ledtråd på ostronet . 
Är det inte på havets botten ? 
Jo , men jag har kanske hittat nån som känner havet . 
Zappos då ? - Undantaget . - Hon är här . Jag måste gå . Hejdå . 
Hej . 
Förlåt att jag inte hälsade på dig ... Förlåt , jag heter Julio . 
Hej , Deedra . Trevligt att träffas . Tack för att du tog fallet . 
Javisst . Bryce ! - Var fan är han ? - Förlåt ! 
Jag har ditt vatten . 
- Mitt vad då ? - Ditt vatten . 
- Du bad om vatten ? 
- Jag var sarkastisk , Bryce . 
- Tycker du inte om mitt skämt ? 
- Jo , det gör jag . Det verkar inte så . 
- Sak samma . Okej , Julio . - Ja . Du tappade ett örhänge i havet . Ja , det gjorde jag . - Det är ungefär tre centimeter . 
- Får jag se bilden ? 
Jag skulle mejla dig igår om det . 
- Visst fick du det ? 
Här . 
Okej , få se här . 
Sen när jobbar fiskar ? 
Borgmästaren sa att om folk förväntas hålla vattendragen rena , så borde fiskar och annat vattenfolk dra sitt strå till stacken . 
Okej , Bryce . - Bryce ! 
- Förlåt , jag är här . 
Örhänget är tre centimeter . Guld . 
- Skriver du ner det här ? - Ja . 
Ja , det gör jag . 
- Format som ett ostron . - Japp . - Med diamanter . 
- Japp . - Har du en extra penna ? - Bryce ! 
Ungefär hur många ? 
Är det viktigt ? 
Varför inte ? 
Jag vet inte . Förlåt . Okej . 
Diamanter . Flera . 
- Och en pärla . 
- Japp . Pärla . Jag ska komma ihåg det . Okej . Vi hör av oss när vi hittat det . 
Bryce , nu går vi . 
Deedra sviker dig inte . 
Jag bara undrade , vad vill du ha till lunch ? Jag vet inte . Kanske fisk ? 
- Julio ? - Ja ? De har stängt av varmvattnet . 
Och varför letar du efter ostronet ? 
De snälla människorna på Zappos ska fixa ett undantag åt dig . 
Det kan ta flera månader . 
Bibo kan inte ta det här nu . Bibo har en viktig provspelning . 
Nästa L-tåg anländer om 178 minuter . 
Vad ska du göra idag , raring ? 
Jag vet inte . 
Du kanske kan söka jobb . 
Ofattbart att den där supermänniskan inte gav dig tillbaka jobbet på köpcentret . 
Du behöver Gud . 
Följ med mig till kyrkan . 
Jag tror inte på sånt . Förlåt . 
Jag är inte sugen på nåt . 
Varför går du inte till Central Park . Det är fint . 
Det är inte Florida men ... New York är inte så illa . 
När jag bygger ett sandslott , hoppas jag att det är kvar nästa år . 
Visst är det kul ? 
Vet ni vad som är skrämmande ? Jag går redan i terapi . 
Jag är yngst och behöver inte bevisa det . 
Älskling , du är inte så ung . 
Inse det . Det är lättare att hata mig än dig själv . 
Varför säger du det inte rakt ut ? 
Jag anlände till Biancas restauranginvigning ... 
- Dina ! - Hej , Bianca . 
... lagom sent . Och jag blev väldigt störd av vad jag såg . 
Bianca . En fråga . Vad har Genevieve för planer för det där hörnet ? 
Vilket hörn ? 
Hörnet därborta . Det är tomt utrymme . Vad är tanken bakom det ? 
Folk förväntas äta här . Hålet kommer att störa dem . 
Kan jag hjälpa dig , Dina ? 
Du behöver inte bli så uppjagad . Jag ställde bara en fråga . 
Jag designade Biancas restaurang . 
Jag vet nog vad jag gör . Jag gick på SCAD . 
På nätet . 
Bombnedslag . 
Utbildningen var på nätet , men datorn var ... stor . 
Tjejer , snälla . Det är en viktig kväll . Kom igen . 
Så för att glömma allt drama i stan tog jag med tjejerna till Sandcastles villor och golfklubb på Bahamas för en liten tjejresa . 
Förhoppningsvis stannar allt drama kring hålet , kvar i New York . 
Jag packade min bikini , min solhatt och allt drama kring hålet . 
Visst är det kul ? 
Det är fantastiskt . 
Och se , Genevieve , alla hörn är fulla . 
Det verkar som att allt drama kring hålet inte stannade i New York . 
Jag pratade inte om det . Du pratar om det just nu . 
Jag säger inte ett ord , raring . Allt är i ditt huvud . 
Prata inte med mig när du pratar med mig . 
Donnie ... ge dem mer champagne . 
De är redan rätt så fulla , sir . 
Herregud , är de ? 
Frågade jag det ? 
Duktig pojke . 
- Du behöver inte bli uppjagad . 
- Det är jag inte . - Du bara skapar drama . 
- Nåväl , Genevieve . Jag har funderat . Det är rätt sjukt att jag tog en chans på dig . 
Alla blev störda av hålet . 
Vad är det som pågår ? 
Låt oss avsluta för dagen . 
Hon är galen . 
Jag designade en vacker restaurang åt henne . 
Tjejer ... Mitt kreditkort har ingen gräns . 
- Säg inget . - Vad är det här ? 
Vem är jag ? 
Allt kommer att bli bra , men du måste hålla dig lugn . 
Stänger av strömmen . 
Jag stannar och stänger . 
- Lyssna , Genevieve . - Vad då ? Allt är okej . 
De ser oss inte . 
Kamerorna är avstängda , men du måste hålla dig lugn . Skrik inte . 
Glen , det är jag . Riktiga Bianca . Andas bara . - Javisst . - Andas bara . Genevieve , du måste se det här . 
Åh , Gud . Om du ser det här är jag så ledsen . 
Jag gjorde mitt bästa men jag misslyckades . Och ... eftersom du ser den här videon betyder det att du inte längre är under deras kontroll . - Hans kontroll . - Vems då ? Hur ? 
Jared , producenten . 
Du har varit fast i hans sjuka lilla pjäs . 
Ditt liv har varit en simulation . 
Men nu är ni två vakna . Jag kan rädda er . Vi kan fly . 
Du verkar bekant . 
Vad heter du ? 
Brandon . 
Mina damer , imorgon händer det . Jag kommer att ha kontroll över dörren . Jag byter ut koden och lämnar dörren olåst . 
Allt ni behöver göra är att ta er igenom en dag till , okej ? 
Vad ni än gör , gå inte in i Jareds kontor . 
Jag är så glad att jag bokade Benihana-upplevelsen för att komma bort från allt drama i stan . 
Jag är dålig i magen . 
Jag sa ju , Rellany . Jag kan inte äta " tortellias " . 
- Var är Brandon ? 
- Övervåningen , med chefen . 
Jag undrar vad han gjorde ? 
Genevieve , du brinner ! 
Din hand ! 
- Hämta lite vatten ! 
- Jag har inte vatten . 
Nån har druckit lite för mycket . 
Stänger av strömmen . 
Snabbt ! 
Det är olåst . - Det är olåst . Kom så går vi . 
- Vänta , jag måste försöka . 
Vi har redan försökt . Nu går vi ! Gen ! 
Nej . Inte utan Brandon . 
Han hjälpte oss . 
- Gen ! - Jag lämnar inte honom . 
Brandon ? 
Var är Brandon ? Var är Brandon ? 
Gud , du är så dum . 
Ja och nej . 
Det är jag , Genevieve . Din skapare . 
Din Gud . 
- Gen ! - Vad ? 
Vad är det här ? 
Hej , Bianca . 
Du ser fin ut . Vad ? Vad är det som pågår ? 
- Varför verkar du så bekant ? 
- Visst gör jag det ? 
Kanske för att ni alla har lite av källkoden i er . 
Källkoden ? 
Ja . Källkoden . 
Den ursprungliga , sanna , rika kvinnan från New York . 
Vacker . Elak . Min mamma . 
Människohjärnan är ... en otrolig sak . 
Man kan utvinna hela världar även efter att kroppen är borta . 
Jag utvinner hennes hjärna för era beteendemönster . 
Det är lätt att hitta en elak , rik dam , men för att skapa en mamma , en mor , så måste jag gå direkt till källan . 
Era hjärnor är sammanflätade med hennes . 
- Ser man på , det är Kycklingben . 
- Kalla mig inte för det , mamma ! Okej ? 
Du vet att det är genetiskt . Du vet att jag fick dem från pappa . Det är inte mitt fel att ni hatar varandra . 
Din mamma brukade låtsas vara sjuk på din födelsedag så att hon fick all uppmärksamhet . 
Hon låtsades vara gay när du kom ut . 
Det räcker ! 
Det räcker , okej ? 
Inget av det spelar nån roll längre eftersom nu ... får jag leka med henne genom er för alltid . 
- Vi går . - Gå ? 
Är det vad du vill ? Ja . 
Jag menar ... Okej . - Dörren är därborta . 
- Gudskelov . 
Jösses . 
Ha så kul i fängelset . 
Glömde ni ? 
Ni är här för att ni skrev på ett kontrakt . Minns ni ? 
Visst är det här bättre än att hamna i fängelset för skattebedrägeri ? 
Mina damer , var inte rädda . Jag och Onkel Sam har en överenskommelse . 
Ni är ju trots allt ... vår största export . En åtråvärd livsstil . 
Men varför befriade du oss ? 
Varför gör du det här ? 
Ibland är det bra att skaka om buren . 
Ert försök till frihet var den perfekta säsongsfinalen . 
I varje fall , vad tycker vi ? 
Några fler säsonger ? 
De har nog inga fodralklänningar i häktet . 
Härnäst på The True Women of New York . 
Igår kväll tänkte jag på min barndom , och jag minns inget . 
Jag mindes inte ... mina föräldrar . 
Nu börjar hon igen . 
Jag tycker att det är smaklöst att inte färga hårrötterna inför en utekväll . 
Det här kallas för en look . 
Förlåt . 
Så de väckte honom med avsikt ? 
Det var som ... en cirkus . Jag älskade det ! 
Så ... berätta hur det känns att äntligen se dig representerad och ... gör mig en tjänst . Säg nåt på spanska . 
Det känns otroligt att äntligen få ett manus som representerar mig . 
När jag fick det så sa jag : " Ay dios mío . " 
Julio , vill du visa henne hur vi egentligen föreställer oss repliken ? 
Abuela , jag gömde mig inte i skafferiet . 
Det måste vara mer som i Pixars animerade filmer , typ ... 
Abuela , jag gömde mig inte i skafferiet , jag letade efter ... salt ? 
Stämmer det att dina tamales skapades med magi ? 
Utsökt . 
Hon är rätt för rollen . 
Adios . 
Vi låter bli att göra den här showen . 
Jag har andra manus . 
Minns du delfinen som fastnade i Gowanus-kanalen i södra Brooklyn ? 
Det skulle vara en riktig bra film . En tre timmar lång film . 
Ingen vet hur delfinen kom dit . 
Okej , förlåt . Lägg av . Sluta . 
Det kommer en tid då du måste växa upp och sälja produkter . Det var otroligt . Vilken förvandling . 
Jag såg dig genom glaset . 
Hur ser din process ut ? 
Jag studerar människor och sminkar . 
Så fantastiskt . 
Jag älskar att prata med skådespelare och lära känna dem . 
Självklart så fick du rollen . 
Ja , det stämmer . 
Jag behöver se ditt filmfack-kort och bevis på existens . 
- Jag har inget sånt . - Vad ? 
Jag är en robot . 
Jag försökte ansöka , men blanketterna har ingen ruta för Bibo . 
Ni vill ha mina idéer , men ni vill att de passar in i er mall . Så det finns inget utrymme för nåt nytt . 
Bibo ? 
Vad är det som pågår ? 
Ett oanvänt Zappo-manus ? 
AVVISAD " Avvisad . " " Kasserad . " " Inte en intressant historia . " 
Bokstaven Q ? " Lejonkungen ur en zebras synvinkel ? " 
MISS VANESJA FRÅGOR ? RING VANESJA OCH FRÅGA EFTER VANESJA Taxi . 
- Vad ? - Ja . 
Jag heter Carl och ringer från Carls telefon . 
Jag hittade ett manus skrivet av en " Julio " ? 
Jag lyssnar . 
Jag ser mig själv i dessa historier och tror att andra som jag skulle hålla med . 
Vi kan nog komma på nåt . 
Så löjligt . 
Han provspelade för rollen . Han fick rollen . Du gillade honom . Ge honom rollen . Jag har en idé . 
Vi kan inte anlita honom som skådespelare , men vi kan anlita honom som rekvisita . 
Så förolämpande . Bibo går inte med på det . - Överenskommet ! 
- Bibo ! Så galet . Jag gör det här utan bevis . Varför kan inte Bibo ? 
Ditt bevis-ärende är under behandling . 
Vi kan säkert hitta ett undantag . 
Bibo vill inte vara ett undantag . 
Bibo vill vara en skådespelare . 
Inkommande samtal . 
En sekund . Ja , hej . Hallå ? Ett ögonblick , tack . Nej , vänta . Det är Julio . Gäller det mitt labbresultat ? 
- Jag sa ett ögonblick tack . 
- Sätter du mig i telefonkön ? - Det var du som ringde ... - Åh , herregud . Jag hatar dem . Hörde du att Nautica var " sjuk " idag . 
Den subban är inte sjuk . 
- Ja , hon har nog bara fått flatlöss . - Ja . 
Vad är det för lukt ? 
Det är nog ett oljeutsläpp . 
Jag tänker inte dö av ett oljeutsläpp som mina föräldrar . 
Jag är så ledsen . Du förtjänade inte det . 
Rättsväsendet log inte mot oss idag . Men jag tycker att vi tog ett litet framsteg genom att belysa ... orättvisor ... 
BEVIS PÅ EXISTENS Vilken osis . 
Jag fattar att Dodo var vresig , men kom igen . Nåväl , nu får nissarna en julbonus . 
De fick inte det förut , så alltid nåt . 
Glaset är halvfullt . Vilken optimist du är , älskling . - Jag älskar det . - Ja . Förlåt . Hej , älskling . Välkommen till Chesters . - Gör du leveranser idag ? - Ja . Tack . 
Okej , oroa dig inte . 
- Chester ... - Vad ? ... det står inget pris i appen . 
Hur mycket kostar det ? Nej , raring . Det är mitt företag . Jag bestämmer . 
Och idag så ger jag dig lite rabatt . 
Okej , bueno . 
Ge mig några nachos . - Jag är hungrig . - Kan jag också få nachos ? 
Vi beställer en till . Hej . Förlåt . För Carl . Jag är Carl . Ja , Carl . Jag vet . Därför är jag här . 
Chester , jag är två timmar försenad . 
Se på dem . Så små och patetiska . 
Dustin , älskling . Jag måste erkänna en sak . 
Den viktiga presskonferensen , jag ... - Jag vet inte vad den handlar om . 
- Ingen fara . 
Jag har en stor idé . Jag har tänkt på den hela morgonen . 
Japp . 
Du vet min roll som en hemlös , gay tonåring i Fittiga Rikemansbarn : Magiskolan ? 
Ja , såklart . 
Det känns fel . 
Jag blir superrik genom att exploatera mindre lyckligt lottade personers svåra belägenhet . 
Älskling , vem lärde dig " belägenhet " ? 
Och alla firar mig . 
Skit i det . 
Jag får betalt . 
Och tv-bolaget , det jävla tv-bolaget tjänar pengar på det . 
De stora oljeföretagen köpte tv-bolaget . Publiken som ser showen tänker : " Oj , hurra ! Vi ser framsteg . " 
Men de inser inte att när de ser på showen så ökar de välståndsklyftan genom att berika just de personer som förtrycker dem som de påstår sig företräda . 
Visste du inte det ? 
Här är min idé . 
Tänk om vi slutar göra showen tills folket i toppen lovar att omfördela vad de tjänar ? 
Vi kan rada upp oss , gå arm i arm , hålla en riktig " bojkitt " . 
- En vad då ? 
- Jag kan få med mig hela ensemblen . Vi kanske kan lyckas få hela branschen att betala alla lika . 
Dustin , älskling . Jag är så stolt över dig . 
Låt oss offentliggöra det . 
- Jag hittade ostronet . 
- Åh , Gud . Jag är på väg för att göra ingreppet . 
Nästa gång du ser mig , har jag ingen kropp . 
Gör inte det . Läste du artikeln jag skickade dig - om de platserna ? - Nej ? Rubriken säger att de utvinner dina färdigheter för att skapa programvaror till att byta ut folk . Gör inget dumt . 
Jag måste gå . Ciao . 
Okej , precis som vi övade det . Från hjärtat . 
Ja . Okej . Uppfattat . 
Tagning . 
Yo , läget , era dammiga puckon ? 
Jag har nåt stort att berätta för er idag . 
Det blir helsjukt . 
Säg inte puckon . 
Okej , jag kan göra det . 
Innan vi gör det här , kan vi bestämma semesterdagar ? 
Jag vill köpa den där villan i Toscana . Jag vill inte förlora den . 
Jag vet inget om nån villa . Vad då ? Varför inte ? 
Med den nya omfördelningen av pengar så kommer du inte att ha - en massa pengar liggandes . - Vänta lite . Blir jag typ pank ? 
Nej . 
Nej . 
Du kommer att ha tillräckligt . Du kommer att åka på semester och vi kommer ... att hitta ett hus till dig . Men ... inte en villa . 
Inte en villa ... 
Och många gåvor . Du kommer att få många gåvor . 
Som den här . Den kom med posten idag . 
Den är nog från en kvinnlig beundrare . 
Ja , antagligen . 
Okej . Låt oss sätta igång med presskonferensen . 
Jag är så stolt . Du ger mig ett syfte . 
Dustin ? 
Blås av den . 
Presskonferensen . Skit i den . 
Varför det ? 
För att ... DU FÖRSÖKTE OCH DET RÄCKER . Jag försökte . Och det räcker . 
Gör det ont ? 
Vill du svara innan du blir av med fingrarna ? 
Hallå ? 
Det passar inte nu . 
- Jag håller på att laddas upp . 
- Är det mr Julio Torres ? 
Jag ringer från Direkt-läkare angående dina resultat . 
Allt ser bra ut . 
- Ursäkta , vad sa du ? 
- Allt ser bra ut . 
- Ursäkta , vad sa du ? 
- Ja , den är godartad . Ha en bra dag . 
Hej . Så det här är inte den saknade delen . 
- Vad menar du ? 
- Den är inte en del av antikviteten . 
Är du säker på att det här är ostronet du letade efter ? 
Ja . Jag är säker . De kollade mina fingeravtryck . 
Okej , ja , den här är från Amazon . 
Så den är inte unik . 
Okej , låt oss börja med att riva ner stället . 
Bibo ? Är du här ? 
Är du hungrig ? 
Jag och Vanesja har en middagsträff för att diskutera mina idéer kring vattenfallen . 
Ett av dem rinner i sidled . 
Bibo ? 
Bibo ? TVÅ MÅNADER SENARE Gjorde du Hur jag kom ut för min Abuela ? - Ja . - Vilken fantastisk show . 
Jag har inte sett den . 
Men bra att du har beviset , speciellt nu då du behöver det för att ... typ rösta och sånt . 
Japp , jag fick precis ett kreditkort och lade till Netflix på det . Häftigt . Du är officiellt hyresgäst ... BEVIS NUMMER 27-44678 NAMN : JULIO TORRES ... av enhet 72 . 
Hem ljuva casa . 
Känn dig som hemma . 
- Hej . - Hej , min lilla stjärna . 
Jag har en överraskning till dig . Jag hittade några människor som gillar dina idéer . 
Kom till lågstadieskolan och träffa dina nya medarbetare . 
Jag är bara före min tid . Tarmflora . 
Du är sen . 
- Till vad då ? 
- Din show . 
Jag måste vara längre bak i alfabetet . 
Sak samma , knäppis . 
Är det inte tjejen som dödade killen i badrummet ? 
SMÅ PJÄSER AV JULIO Kay gör samma sak som du . Du och din patetiska pinne . 
Macro , vakna . Stäng av teven . 
Jag har fått syn på Bibo . 
Bibo flyger in . Och Bibo har landat . Uppfattat ? Bibo har landat . Du måste säga uppfattat . Uppfattat ? 
Edwin ! Den stannar inte på mitt lilla huvud . 
Ingen fara . Oroa dig inte . - Jag fixar det . - Älskling , hur ser jag ut ? Vacker . 
Har Bibo två roller ? 
Föredrar Carl honom ? 
- Jag spelar bara en roll . 
- Nej , bebé . Fokusera inte på Bibo . Fokusera inte på nån annan . Fokusera på dig själv . 
Ja . Tack . 
Har du ätit ? - Ta en av mina energikakor . - Okej . 
Lycka till . 
- Hur lång är den ? - Den borde ta slut ... nu . 
Släng allt skräp ni har . 
Ingen återvinning i byggnaden , tack . 
- Tack . - Mycket vackert . - Mycket vackert . - Ska vi ... Ja , kom så går vi . - Hejdå . - Hejdå . Ciao . 
Jäklar . Jag måste hämta min mobilladdare . 
- Vi ses ute . - Okej . 
Hej , du . Skrev du det här ? 
- Ja . - Varför ? 
Bad du ens om tillåtelse ? 
Varför är du klädd så ? 
Det är oacceptabelt . Boka flyget . 
Ja . Hej , Vanesja . 
Jag måste ringa dig tillbaka . 
Varför följer du efter mig ? 
Du gav en otrolig föreställning . Vanesja . 
Jag frågar dig en gång till . Varför följer du efter mig ? 
Jag var branschens bästa agent ... tills min lata artist-syster började göra en föreställning om mig och stal mitt liv . 
Bibo ? 
Vanesja . 
Du är bra . 
Bibo är också en artist . Jag har också idéer . Jag gör bara andra grejer hela tiden . 
Jag är med i fotbollslaget , så jag ... Jag förstår . 
Här . Ta mitt läkarintyg . Du är befriad . 
Visa dem det . Gör inget du inte vill göra . 
