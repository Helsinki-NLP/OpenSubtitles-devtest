- Två till . 
- Ska bli . 
Bucky har då all tur . 
Ja , hon är snygg . 
Jag menar inte det . Den tursamma fan åker imorgon . 
Han blir bara ett stenkast från tyskarna medan vi andra harvar på med övningsuppdrag över Nebraska . Oroa dig inte . Vi är snart där borta och fäller bomber . - Ja . - Bucky , vi bjuder på nästa omgång . 
Han har aldrig bjudit förut . 
Så du kallas Bucky och han Buck ? 
Det är en lång historia . 
Visst är de ett fint par ? Jag borde ha presenterat dem tidigare . 
Han åker imorgon . 
Alla behöver nån att skriva till där hemma . 
Jag vet inte om John Egan är brevskrivartypen . 
Om han träffade en flicka som är värd att skriva till , så kanske . 
En flicka värd att skriva till är svår att hitta . 
Inte om man letar på rätt ställe . 
Jag förstår vad du menar . 
Så skriver du till mig ? 
Det är redan gjort . 
Har du skrivit till mig ? Ja . Vad står det i brevet ? 
Tja , du får vänta och se . 
När får jag brevet ? 
När jag skeppas iväg . Kanske om två , tre veckor . 
Jag ska sakna dig varje sekund . 
Okej . Mina herrar , en skål . 
Buck , Marge ... hallå , turturduvor ... vi skålar för Bucky här borta . 
- För vår nya trådjaktledare , Bucky . - Skål . Okej , major . Befäl för alla fyllon i 100:e . 
Nån måste ju göra allt i ordning för er andra träskallar . 
- Skål , major . - För 100:e . 
- Ja , för 100:e . - Lycka till , sir . - Tack . - Spara några tyskar åt oss . 
Vi går till Slooter . Hänger ni med ? 
Nej , jag måste flyga tidigt . - Buck ? 
- Jag tror inte det , killar . 
Vi ses imorgon då . Hej då , Marge . 
Bucky , vi ses i England . 
Kom ihåg att jag vill ha extra filtar och en brits med utsikt . 
Det ska vi fixa . 
Han vägrar berätta om smeknamnen . 
Berätta nu , Marge . 
- Ska jag ? - Visst . - Okej . - En lång historia , som sagt . 
De träffades under grundutbildningen innan kriget började . 
John har kallats Bucky sen han var barn . 
- Visst ? 
- Det stämmer . 
Och Gale ... Tja , Gale har alltid kallats Gale . 
Ända tills ... Första dagen på grundutbildningen kommer en kille fram till mig och säger att jag liknar nån där hemma i Wisconsin som kallas Buck . 
Jag säger att jag heter Gale , Gale Cleven . 
Och ... Men Bucky ger sig inte . Nix . 
Det är " Buck hit " och " Buck dit " . 
" Buck , hjälp mig knyta skorna . " " Buck , hjälp mig flyga det här planet . " 
Innan jag vet ordet av kallar hela jädra 8:e flygflottiljen mig Buck . Så ... Gale är inget vidare bra namn . Vet du vad ? Du borde tacka mig . Jag gjorde dig en tjänst . - Som gav mig samma namn som du ? - Inte exakt samma , och jag rår inte för att du såg ut precis som Buck - från Manitowoc , Wisconsin . - Från Manitowoc . Vem gör så mot sin bästa vän ? 
- Så rart . - Vi behöver musik . 
Okej . Försvinn inte , Gale ... Buck . Du ska dansa med mig innan kvällen är över . 
Tvinga mig inte att dansa , Marge . Välj nån bra låt . 
Artie Shaw , Benny Goodman . 
- Hej . - Det är helt otroligt att vi är vänner . 
Du vill inte dansa med en vacker kvinna . Du varken dricker eller spelar . 
Du gillar inte ens sport . 
Tja , vi är ett av livets stora mysterier . - Den gillar jag . Ja . - Jaha ? Så nu är det dags . 
Det är dags . 
Vi ses om några veckor . Om jag inte hinner dö . 
Tyvärr är du trådjaktledare för 100:e nu . 
Du lär inte flyga uppdrag där borta . 
Alltså , jag pratade med befälhavaren för 389:e , och jag ska flyga med dem tills ni anländer . 
Jag ska vara observationspilot . 
Din jäkel . Tja , nån måste ju känna på lite strid , så jag kan berätta hur det är . 
Våga inte gå och dö innan jag hinner dit . 
Det vet man aldrig . 
Dyk ! Vi måste släcka motorbranden ! 
Kom igen , fortare ! Du måste hjälpa oss ! 
Bra ! Branden är släckt ! Stig ! 
Stig ! 
Stig mer ! 
- Fiendeplan klockan 12 , rakt fram ! 
- Helvete ! 
Vi har mist fjärde vingklaffen . 
Pilot till navigatör . 
Vi måste återvända . Vi behöver en ny bäring ! 
Helvete ! 
Duval här . 
Jag är träffad . 
Jag kommer ner till dig , Duval . 
Bäring rakt västerut . Uppfattat ! Motor två tappar oljetryck ! 
Håll det stadigt medan jag får en ny bäring . 
Andas ! Andas , bara ! Håll ut ! 
- Duval ! Var är du träffad ? 
- Helvete också . 
Håll ut , Duval ! 
Jag är här . 
- Jag kommer inte att klara mig . - Sluta . Du kommer att klara dig . 
Tryck med handen mot såret . Här . Bra . - Okej . - Förstått ? Håll ut , förbanne mig ! 
Hör du det ? 
Se på mig ! Öppna ögonen ! 
Andas , andas ! 
Fiendeplan klockan 12 ! 
Jag fick en ! 
Egan , jag behöver bäringen ! 
Ny bäring : Gira vänster vid 248 . 
Uppfattat ! 
Kom igen . Håll ut . 
- Vi flyger hemåt . - Ja . Ja . 
Fortsätt andas bara ! Det var ett sjujäkla spaningsuppdrag , major . 
Är det jämt så ? 
Undrar du vad du ska säga till mannarna ? 
Säg ingenting . De lär sig . 
Det gör vi allihop . 
100:e bombgruppen sändes till England våren 1943 för att ansluta sig till USA:s 8:e flygflottilj i kampen mot Nazityskland . 
Jag tycker att vi kallar planet Alice From Dallas . 
Alice From Dallas ? 
Det låter inte dumt . 
Alice From Dallas . Alice , vårt palats . 
Visa för major Cleven . 
Lorch , visa majoren . 
Jag vill ha henne tillbaka . 
Sjutusan till kvinna . Hon ger det här planet lite extra muskler . 
KOM TILLBAKA TILL MIG , KEN ! PUSS , ALICE Jag förstår varför du vill döpa planet efter henne . 
- Hon är speciell . 
- Hon är formidabel . 
Amison , är du säker på att vi är i rätt fjord ? 
Absolut . Helt säker . 
Nutting , hur ser det ut bakom oss ? 
Åtta på rad , sir . Uppfattat . 
Få av oss hade varit långt hemifrån , ännu mindre flugit med ett flygplan . 
Vi kom från landets alla hörn , med ett gemensamt mål : att ta kriget till Hitlers tröskel . 
Piloten till besättningen . Vi landar strax i Grönland för lite mat och vila . 
Blondie Tower , Army 233 . En grupp B-17 över Bluie West One . 
Landningsinstruktioner , tack . 
Army 233 , flight Blondie Tower . 
Fortsätt mot landningsbana sex . Klart att landa . 
Klar sikt . Vindar från 330 på 40 knop med vindstötar upp till 50 . 
Höjdmätare 2990 . 
Det är lite blåsigt . Blåsigt ? 
I ' Bama kallar vi det orkan . 
Uppfattat , Blondie Tower . Fortsätter mot landningsbana sex . Klar sikt . 
Vindar från 330 på 40 knop med vindstötar upp till 50 . 
En sjujäkla sidvind . Ökande vindstötar . Var försiktiga . 
Kanske bäst att cirkla runt , major . Välkomna till Grönland . 
Landningsställ nere . Var redo med klaffarna . 
Landningsstället fälls ner . 
Det blir skumpigt . Håll i er , killar . 
Pilot till besättning . Beredskap för landning . 
Vänster nere . Höger nere . 
Sista landningskontroll . Klaffar en fjärdedel ner ? Japp . Klaffar en fjärdedel ner . - Klaffar halvt ner . - Klaffar halvt ner . 
Klart . 
Stig , Veal . Vänd och kom tillbaka . 
BLUIE WEST ONE FLYGFÄLT SÖDRA GRÖNLAND Vår bombgrupp bestod av fyra skvadroner . 
Major Gale Cleven förde befäl över 350:e . 
Han och major Egan var de obestridda ledarna för hela vår bombgrupp . 
Ev Blakely var pilot från Seattle . - Titta här . - Blakely . 
Och generöse Benny DeMarco från Philly . - Major . - DeMarco . 
- En sjujäkla landning . 
- Jag har sett värre . 
- Är det boxningsmatchen ? - Ja . 
- Claytor , du har pengar på den , va ? - Ja . - Men det är dålig mottagning . - Ja , verkligen . 
Dra upp volymen . 
Bombfällarna James Douglass och Howard Hamilton kom från Mellanvästern . 
Hambone . 
- Major . - Japp . Lugn . Jag fixar det . Charles Cruikshank , känd som Crank , var från New England . Tjena , Crank . Ni hade visst en svår landning . 
Min bäste vän Joe " Bubbles " Payne och jag var navigatörer , så lokalisering var viktigt för oss . Major ? Löjtnant Crosby . 
Varifrån är ni ? 
Vi måste sätta en nål i kartan . 
Bubbles och jag ... vi håller traditionen levande . 
- Här är folk från hela landet . - Ja . Casper , Wyoming . 
- Cowboydelstaten , va ? - Japp . 
Tja , ni är visst den förste därifrån , major . Tänka sig . Major . Vad önskas ? 
En vän till mig landade här för några veckor sen . En trådjaktledare . Det skedde visst en incident . 
Är ni vän till Egan ? Major John Egan ? Bucky ? 
Det stämmer , ja . 
Jag vet inte vad han sagt , men jag gjorde inget fel . Nej , han bad mig att ge er den här . 
Som ersättning , sa han . 
Ersättning ? Ja . Och hur skulle den här kunna vara en ersättning ? 
Sergeant , jag vet inte vad som hände , men han sa att den där bör göra er kvitt . 
Titta där . 
Avbruten narvalsbete . Han drog ner den från väggen och lekte enhörning . Han förstörde två soffor och krossade nästan alla glas i baren . 
Jag förstår . 
Jag brukar kunna identifiera en bråkmakare , men din vän verkade okej . 
Tills han började sjunga . 
Ja , det känner jag igen . 
Du behöver inte göra det här . Det är ett fånigt vad . Nu är jag tvungen . Vem ska det bli ? 
- Okej , lugn . - Vem ska det bli ? 
Jag har mött varenda en av er och ni irländare är lika usla på dart som på att slå i en spik . 
Skratta inte . Ni engelsmän är inte mycket bättre . Jack ! 
Men Tommy här är den bästa dartkastaren - i hela East Anglia ! - Du mister ögat . 
Nej då . Jag litar på Tommy . Om han vinner , får jag båda cyklarna . 
Kör i vind , yankee . 
- Båda två . 
- Okej , båda två . 
Och jag får en kyss . Okej , Tommy . Inte mina ögon . Inte mina ögon , okej ? 
Okej , Tommy . När du är redo . Jag har just förlorat två cyklar , Tommy . - Vad är det med dig ? - Tommy ! 
EAST ANGLIA , ENGLAND 8 JUNI 1943 
ENDAST BEHÖRIG PERSONAL - Godkväll , major . 
Är cykeln till salu ? - Inte på några villkor . 
Det var mitt jobb att få kapten Brady och resten av besättningen från Grönland till vår bas vid Thorpe Abbotts i England . 
Men på nåt sätt skildes vi från resten av gruppen bland molnen över Atlanten . 
Svårt nog med obefintlig sikt , men jag hade ännu ett problem : okontrollerbar flygsjuka . Vi har ett elektriskt problem . Vi behöver en bäring . 
Crosby , är du där ? 
Ursäkta . Kan du repetera ? 
Vi har knas på elsystemet . 
Ge oss en riktning medan vi löser det här , Croz . Uppfattat . Avvakta . 
Gira höger till 165 . Kom . Uppfattat . Girar höger till 165 . 
Stänger av det elektriska och startar om det . Vi fixar det här . 
Säkert en av kontrollkretsarna . 
Jag drar ur säkringarna . Det isolerar problemet . Okej . Kör . 
Hur kan du spy än ? 
Din mage måste vara lika tom som vår bränsletank . 
Ja . Ja . - Åh , men för tusan , Croz . 
- Förlåt . 
Jag har spyor över hela mig . Ge mig en trasa . 
- Förlåt , förlåt . - Sätt fart . 
Det stinker . 
Hur går det ? 
Inget elknas såvitt jag kan se . Kanske problem med hjulmotorn . 
Startar om batterier och generatorer . Tillbaka på . 
Varningslamporna av . 
Är det där Englands kust ? 
Crosby , visst är det England ? 
Nej , vi borde inte vara över vatten . 
Sir , vad är bäringen ? 
165 , precis som du sa . 
Men för alla milda makter . 
Fan också . Det är Frankrike ! 
Pilot till besättning , luftvärnseld framför . Håll i er . Fan ! 
Men för fan , Croz . THORPE ABBOTTS FLYGBAS Morris . Tack för cyklarna . 
Jag slår dig nästa gång . Såja . Kom , kossan . 
Här kommer de . Kom , vovven . 
DeMarco ! 
Hej , major . 
Var fick du tag i hunden , Benny ? 
Jag vann honom på tärning . 
Tog du upp vovven över 3 000 meters höjd ? 
Han har syrgasmask . Den kostade mig tre dollar . Men han älskar att flyga . 
- Han ylade hela tiden . 
- För att han är delvis varg . 
Han är en varg som är delvis hund . 
- Vad heter han ? 
- Meatball . 
Välkommen till 100:e , Meatball . 
Kom nu , Meatball . 
Har du saknat mig ? 
Som en sten i skon . 
- Hur har du haft det ? - Hälften av utrustningen har inte kommit . 
Jag fick låna syrgasmasker och fallskärmar av britterna . 
Trådjaktledaren bör sköta det . 
Enligt mig borde de avskeda honom . 
Och vänj dig vid leran . 
Jo , du , har din radiokille hört nåt radioprat från 418:e ? 
Brady saknas . 
Svar nej . 
Jag har en cykel åt dig . 
Behöver jag en cykel ? 
Annars tar det 20 minuter från logementet till mässen . 
Och såna här går inte att få tag i . 
Nu kan du susa förbi ett helt kompani som traskar i regnet på väg till middagen . Du kommer tillbaka och säger : " Tack , Bucky . " 
Räkna inte med det . 
Där kommer Brady . 
Okej , kolla landningsstället . Sänk ner det . 
Uppfattat . 
Vänster ner . 
Bakre ner . 
Men inte det högra . 
Helvete . Höger hjul har fastnat . 
- Blum , veva ner det manuellt . - Ska bli . 
Hafer , hjälp honom . 
Uppfattat , ska bli . 
Ta den . 
Var är veven ? 
Kom igen . Det sitter fast . 
- Kom igen . 
- Jag försöker . 
Ur vägen . Såja . Ge hit den . 
- Har du tag ? - Ja . 
Motorn till landningsstället är paj , eller skruvdomkraften . 
- Är du säker ? 
- Ja , sir . 
Det är helt fast . Det går inte ner . 
Fäll in vänster landningsställ . 
Är du säker ? 
Ja , vi har större chans med en buklandning än om vi landar med ett hjul . 
Clear-up Tower , Army 071 här . Landningsstället fungerar inte . 
Begär landningsinstruktioner . Kom . Uppfattat , Army 071 , klartecken att landa . Räddningsmanskap är redo . Kom . 
Uppfattat , Clear-up . 
Pilot till besättning , var redo för kraschlandning . 
Hörde ni ? Kom igen . Sätt fart . 
247 . Räddningspersonal ... - Okej . Alla ut ! Alla ut ! - Sätt fart ! Alla ut ur planet ! 
- Sätt fart ! 
Fort ! Sätt fart . Spring , annars dör ni . Fort ! - Alla utom fara . - Åh , helvete . 
Enkel sak . 
- Koppla på vajer och bogsera . - Ska bli . Kom . 
Du är navigatör , Crosby . 
Du borde kunna , jag vet inte , hitta England . 
Är alla oskadda ? 
- Ja , sir . - Sir . 
Brady . Kliv in på mitt kontor . 
Hur tappade ni bort de andra ? 
Vi blev skilda åt i molnen . 
Och sen hade vi elfel av nåt slag , så vi försökte få ner landningshjulet i en timme . 
Du vet hur man brukar säga . Det finns två slags piloter , de som har gjort en buklandning , och de som kommer att göra det . 
Major , det ser värre ut än det är . - Okej . Ta hand om det . - Ska bli . 
Du behöver inte urskulda mig . - Det var mitt ansvar . Jag borde ha ... - Det gjorde jag inte . Vi hade ett mekaniskt fel . 
Få bukt med flygsjukan . Eller lämna mitt plan . 
Croz , tog du den natursköna rutten ? 
Nå , tänker du berätta om det där med enhörningen ? 
Enhörningen är min favorit bland utrotade djur . 
Frankrike ? 
- Hur fan bar du dig åt ? - Vad tror du , Bubbles ? 
Jag spydde som en räv . 
Jag trodde att det gick över - när du kom upp i luften . - Ja , vanligen . Men den här gången , med turbulensen ... Jag vet inte . 
Det gick inte över . Jag är säkert den sämsta navigatören i hela flygvapnet . 
Äsch , det finns nog nån som är sämre . - Åtminstone en . - Akta . Fel sida av vägen , löjtnant . - Sir . 
- Välkommen till England . 
De där två har nog sett Test Pilot några gånger för mycket . 
Det har du också gjort . Ja . 
Det hjälpte inte . 
Vi får i alla fall tala om vartåt de ska rikta planet . - Vi ses , Buck . - Tack för skjutsen . Raka vägen i vanliga fall . I ditt fall den natursköna rutten . 
Jaha , den natursköna rutten ? Mycket lustigt . 
Jag borde inte behöva förklara för er det allvarliga i ert ansvar . 
Ni vet att det här inte bara handlar om hur bra er besättning bäddar sängen . 
Det gör jag , sir . 
Därför prioriterar jag flygtimmar framför bäddning . 
Ni har befäl över 35 plan och 350 flygbesättningsmän . 
Pojkar utan stridserfarenhet . 
Deras liv hänger på ordning och disciplin och ert föredöme . 
Ja , sir . 
Med all respekt kunde jag nog vara till större nytta för dem och er som skvadronbefälhavare än som trådjaktledare . 
Att ha en framskjuten position gör en inte till ledare . 
Jag tror helt enkelt inte att jag passar bakom ett skrivbord . 
Jag behöver vara där uppe och hjälpa killarna . 
Överste LeMay har ögonen på oss . Han bara väntar på att få lägga ner 100:e bombgruppen . Det tänker jag inte låta ske . 
Och jag väntar mig att alla officerare ska sätta skuldran till . 
Jag menar er , major Egan . 
Det var allt . Hur är det , sir ? 
Ska jag kalla på doktorn ? 
Det är ingen fara . 
Inom kort väckte de oss för vårt första uppdrag . OFFICERARNAS KVARTER Efter hundratals timmar flygträning i Staterna måste vi tro att vi var redo . 
Vi måste , för nu var det allvar . 
Sir , ni ska flyga idag . 
Major Cleven , sir . 
Det serverades jämt en särskild frukost inför ett uppdrag : ägg , fattiga riddare , pannkakor , en dubbel ranson bacon , färsk grapefruktjuice och några koppar armékaffe . 
Mannarna kallade det den sista måltiden . 
Hoppas att vi alla återvänder helskinnade från ... Chuck , skicka saltet , va ? 
- Oj då . - Jäklar . Han spillde ut saltet . 
Var snäll och kasta saltet över axeln , så vi alla kan fortsätta med frukosten . 
- Vem gjorde det där ? - Jösses . 
- Inte alltihop , Chuck . 
- Det bringar oss inte otur . 
Kasta saltet , sa du . Dumskalle . 
Kasta saltet , sa han . 
- Curt , jag flyger med dig idag . - Här . - Vad sa du ? - Ursäkta , Dick . Då hamnar du i aktern , men du kan ändå skjuta tillbaka . 
- Det är okej . 
- Gör Meatball sig klar ? 
Lemmons eller Wink håller ett öga på honom . 
Följ inte med på det här uppdraget . Ett gott råd . 
Bäst att jag äter några ägg innan alla är slut . 
Gör inte det , Buck . 
De där äggen värptes innan jag kom i målbrottet . Okej , jag hoppar över äggen . 
- God morgon , pojkar . 
- Major Veal . God morgon , sir . 
Har ni sovit gott ? - Jävligt gott . - Som ett barn . 
Flyger nya skvadronsbefälet med oss ? 
Den nya , eller den ännu nyare ? 
Bekymra dig inte om honom . Fokusera på flygningen . 
Jag vill ha så jädra tät formering att inte ett mynt ryms mellan vingspetsarna . 
- Ja , major Veal . - Ja , sir . 
Giv akt . 
Lediga . 
Dagens mål är Bremen . Vi ska bomba ubåtsbaserna vid floden Weser . 
Jag kan inte nog betona det här målets vikt . 
Vi miste nästan 70 fraktfartyg genom ubåtsangrepp förra månaden . 
Och om vi inte kan frakta materiel från USA till Storbritannien , kan vi inte landstiga på kontinenten . 
350:e ligger högst med major Cleven som chefspilot , och 349:e ligger lågt med major Veal som chefspilot . 
Jag är längst fram med löjtnant Dye i 351:a . 
Efter formationen följer 100:e med 94:e , 95:e och 96:e bombgruppen . 
Vi flyger lägst . Och längst bak . 
Det blir en total flygstyrka på 78 tunga bombplan . 
- Helvete . - Major Bowman , vår underrättelseofficer , fortsätter genomgången . Och kapten Becker avslutar med väderutsikterna . Major . 
Tack , sir . 
Lyse , tack . 
Notera luftvärnspositioner både till sjöss och på land längs Frisiska öarna , från Norderney till Langeoog . 
Över fastlandet kan vi vänta oss kraftig luftvärnseld från Wilhelmshaven , hela vägen till Bremen . 
Identifierade batterier utgörs av 88 och 105 mm-kanoner vägledda av Würzburg-radar , så de lär spåra er . 
Navigatörer , bombfällare , när vi är klara här , rapportera till högkvarteret för särskild genomgång . 
Alltså , er referenspunkt är den nordvästra delen av Bremen , här . 
Målkarta , tack . 
Från den referenspunkten är det raka vägen 15 km till målet . 
Det här är dockorna på östra sidan av floden . 
Den här centrala dockan är ert huvudmål . 
Er bäring fram till inledningen är 218 grader . 
Direkt efter vändningen följer ni floden . 
- Varsågod , major . 
- Tack . 
Få höra , Curt . Vad är dagens citat ? 
Jag ska flyga som en ängel idag , inte dö som en . Major , den är för trång . Jag får inte på mig den . 
Buck , hjälp mig med jackan . Jadå . 
Jag gillar ditt rakvatten . 
Bra . Så här nära mig vill jag att du flyger idag . 
- Precis som vi har övat . 
- Ja , sir . 
God morgon , mina herrar . 
För er som inte känner mig , är jag fader Teska . 
Mitt kontor är strax intill . Kapten Phillips också , ifall nån behöver oss . 
Tack , pastorn . Det ska vi komma ihåg . 
Buck . 
- Hej . - Allt väl ? 
Vad är det här ? Gör du upp gamla räkningar ? 
Det är min tursedel . Din tur ... 
- Jösses , John . 
- Här . Ta den . 
Jag har haft den med på två uppdrag . Allt har gått bra . 
Titta , två hörn avbitna , ett för varje uppdrag . Här är jag , oskadd . Ta den . 
För god tur . 
Okej . Vi ses sen . 
- Okej . - Vi ses sen , allihop . 
Jag ska upp dit . 
Samlas kring mig . 
Som ni vet är det vårt första uppdrag här . 
Jag litar på att ni minns er utbildning och kan era uppgifter . 
Nu ser vi till att klara uppdraget och fälla bomber på nazistskitarna , så får vi åka hem tidigt . 
Ja , sir ! 
Majoren här ska flyga med oss . Major ? 
Första gången det är allvar , pojkar . 
Vi radar upp målen och mosar dem . 
Ja , sir . 
Okej . Så varför står vi kvar här ? 
- Allt okej här bak , Dickie ? 
- Skojar du ? 
Lika bekvämt som en svit på Ritz . 
Tack . - Mina herrar . 
- Sir . En välsignelse att ha er ombord , sir , Jag förnimmer Guds ande i er . 
Ja , i oss allihop , kompis . 
Du höll sätet åt mig . Ja . 
Hellre det än att ha dig sittande i mitt knä tills jag flyttar mig . 
Redo för checklistan . 
Form 1A ? 
Klart . 
Bränsleventiler och brytare ? 
Båda bränsleventiler och brytare i avstängt läge . 
Mellankylarna kalla . 
Gyro ? 
Brytare för bränsleavstängning ? 
Alla fyra öppna . 
Kylklaffar ? 
Öppna vänster och låsta . 
- Reglageställ ? - Reglageställ stängda . 
Huvudströmbrytare och tändlås ? 
Batterier på . Klart . 
Hjälppumpar , tryck ? 
Pumparna på . 
Bränslemängd , bra . 
Okej , löjtnant , redo att starta motorerna ? 
Ja , sir . 
Starta ettan . 
Fint att ha er med , överste . - Starta tvåan . - Startar tvåan . 
Bränsletryck , oljetryck ser bra ut . 
Starta trean . 
En B-17 hade 12 maskingevär som skydd åt alla håll . 
Vi kallade dem Flygande fästningar . 
Men nyckeln till att överleva var att flyga tätt och kunna ge försvarseld från en tät formation . 
Det var viktigt , för om vi skingrades kunde de tyska stridsplanen skjuta ner oss ett i taget . 
Ge dem vad de tål ! Ge grönt ljus . 
Då kör vi , pojkar . Sextio . 
Nittio . 
100 . 110 . 
Okej , pojkar . Nu kör vi . Fyrtio . Femtio . 
Sextio . Nittio . 100 , 110 . 
Vi stiger än , pojkar . Tre timmars färd till målet . 
Checklista efter start . 
Stigeffekt inställd . 
Kylklaffar okej . 
Höger landningsställ uppe . 
Vänster landningsställ uppe . 
Bakre hjulet uppe . 
Okej , Bosser , dags att klättra ner . 
Okej , Curt , jag har kontroll . 
Pilot till besättning . Tretusen meter . 
Syrgasmasker på och rapportera . 
Kulsprutetornet , klart . 
Akterskytten , klart . 
Midjeskytt höger , klart . 
Midjeskytt vänster , klart . 
Radion , klart . 
Flygmekaniker , klart . 
Navigatören , klart . 
Bombfällaren , klart . 
Best , skjut av en lysraket . 
Få se om vi kan komma i formation i den här ärtsoppan . 
Ska bli . 
Är det där en lysraket ? 
Nosen till besättning , jag såg en lysraket rakt under oss . 
Uppfattat . Såg du från vem ? Svar nej . Rena ärtsoppan där ute . 
Jösses ! B-17 rakt fram lågt . Rakt under oss . 
Roy , stig ! 
Jäklar ! En Flygande fästning strax ovanför oss . 
Uppfattat . Jag ser den . 
Akterskytt , rapportera . Men för tusan , går vi fria ? 
Akterskytt till pilot , vi går fria . 
- Det var nära ögat . 
- Det där är Clevens plan . 
Jag känner igen lukten av rakvattnet . Skojar du ? 
Du sa ju åt honom att flyga nära . 
Inte så nära . 
Pilot till besättning , vi har en timmes färd kvar i den här ärtsoppan . 
Håll korpgluggarna öppna . 
Jösses . Vi måste hinna ifatt resten av gruppen . Vi är långt bakom . Formationen är en enda röra . Motor ett går orent . 
- Den stannar . - Helvete . 
Pilot till akterskytt . Vad kan du se bakom oss ? 
Akterskytt till Cleven , från vår grupp har vi sex i formation . 
351:a ligger i formation men 349:e är långt efter . Alla sex . Deras etta , Veal , verkar ha problem . 
Uppfattat . Redmeat Etta , Surface Etta här . 
Vad pågår där bak , Veal ? 
Surface Etta , vi har motorproblem . Jobbar på det . Uppfattat . Du måste ta ett beslut , Veal . 
Du utsätter din skvadron för fara . 
Pacer Etta , uppfattat . Sir , vi ligger långt efter gruppen . 
Ju längre vi väntar , desto längre tar det för dem att hinna ikapp . 
Fan också . Stäng av den . 
Stänger av bränslet . 
Pacer Etta , Redmeat Etta här . 
Vi har mist motor ett . 
Vi kan inte hålla farten . Vi återvänder hemåt . 
Uppfattat , Surface Etta . 
Redmeat Två , vi har motorfel . Jag återvänder hem . Du är gruppchef . 
Uppfattat , ska bli . 
Pilot till besättning , vi intar ledarposition för Redmeat . 
Gå till maximal motorkraft . 
Övervaka vår förbrukning . Det tar mycket bränsle att komma ikapp resten av gruppen . - Eld ! - Eld ! 
Var beredda . Inkommande luftvärnseld . Håll i er , pojkar . 
Kanontornet till besättningen , luftvärnseld klockan elva lågt . 
Luftvärnseld klockan tio högt . Klockan fyra högt . 
Luftvärnseld överallt . 
Må Gud näpsa honom , ber vi ödmjukt . 
Och må du , fursten över den himmelska härskaran , med Guds kraft , kasta Satan ner i helvetet . 
Navigatör , hur lång tid till målet ? 
Cirka elva minuter . 
- Uppfattat . - Elva minuter ? 
... den himmelska härskaran , och alla onda andar ... Jävlar ! 
... som drar runt på jorden och försöker snärja själar . Amen . Helvete . 
Bombfällare till befälspilot , vi bör vara över målet , men jag ser inte ett jäkla dugg . Ska jag fälla ? 
Det går inte . Det går inte . - Sir ? - Jag vägrar fälla bomberna om vi inte kan se det jäkla målet . 
Navigatör , hur verkar det sekundära målet ? 
Navigatör till befälspilot , samma läge . 
Sikten är noll , sir . 
Befälspilot till besättning , jag avbryter uppdraget . 
- Navigatör , förbered ny bäring . - Uppfattat . 
Zootsuit Etta till Zootsuit Två . 
Roger . Uncle . Fox . Xray . Upprepar . Roger . Uncle . Fox . Xray . - Fan också , befälhavaren avbryter . - Helvete ! 
Surface Etta till Pacer Etta , uppfattat . 
Pilot till besättning , uppdraget inställt . Upprepar , uppdraget inställt . Luftvärnselden har slutat . 
Ni vet vad det betyder , pojkar . Okej . 
Var redo , killar . 
Uppfattat , major . 
Befälspilot till akterskytt , vad ser du bakom oss ? 
Jag ser inte 349:e . De är fortfarande långt efter . 
Clevens grupp ligger tätt med oss . 
Uppfattat . Håll ögonen öppna efter fiendeplan . 
När som helst nu , pojkar . Håll korpgluggarna öppna . 
Övre kanontorn till besättning , klockan tolv högt . 
Jösses , vad snabba de är . 
De ger sig på Veals grupp . 
Jaktplan , klockan tolv högt ! 
Helvete . 
Adams , hoppa . Ser nån några fallskärmar ? 
Akterskytt till pilot , jag ser inga fallskärmar . 
Uppfattat . Fortsätt varna för jaktplan . 
Jaktplan ! Klockan tolv högt ! 
Schmalenbach är träffad . Gode Gud . Schmalenbach störtar . 
Jävlar . De kommer rakt mot oss . Jösses . Mullins . Cleven till akterskytt , vad ser du bakom oss ? 
Akterskytt till Cleven , 349:e är i en molnbank . 
Jag kan inte se dem , sir . 
Fiendeplan kommer mot oss . 
Jaktplan klockan sex . Klockan åtta ! 
Fan också . Den kärvar . 
Helvete ! 
Kom igen ! Kom igen ! 
Fan också ! Jösses . 
Akterskytt , rapportera , Dickie . 
Akterskytt till Cleven , jaktplanen är borta . 
Jag ser bara två kvar från 349:e , sir . Tre plan har skjutits ner . 
Dickie , upprepa . 
Det är bara två kvar från 349:e , sir . 
Jösses . 
Kulsprutetorn till pilot . Sir , de sköt hål i tornet . Jag fryser ihjäl . Kan nån få mig upp härifrån ? 
Killar , hjälp Bosser upp och få honom varm . 
Hur är det med Bosser ? 
Vi jobbar med honom , sir . 
Din dräkt är sönderskjuten . Klart att du fryser . 
Ge honom en filt . 
Håll ut , pojkar . Vi återvänder till basen när vi har dumpat bomberna i Kanalen . 
Ingen motorkraft , och så gav den upp helt . 
Verkligen otur på första uppdraget , major . 
Länken till förgasarblandningen fick ett tändstift att sota igen . 
Det tar bara några timmar att laga . 
Sju , åtta , nio , tio , elva , tolv , tretton , fjorton , femton . 
- Vi hjälper dig . - Sätt fart . 
Helvete . Överste ? 
Överste , hur är det ? 
Jösses . Hur är det , sir ? 
Befälhavaren behöver hjälp ! 
Det kommer inga fler . 
- Jag räknar till 15 . 
- Jag med . 
Nitton lyfte , ett avbröt . Tre saknade . 
- Alla från Veals skvadron . 
- Kom nu . - Rapporten , sir . 
- Inte nu . 
Okej . Upp på lastbilen , för fan . Van Noy ! Hallå ! Glen ! Glen ! 
Hallå , Veal . Lugna ner dig . 
Alla håller tyst . Upp på lastbilen . 
Inte ett ord till . Spara det till utfrågningen . 
- Van Noy . Upp på lastbilen . - Till förhöret genast . 
- Inte ett ord till . - Jag vill bara veta - vad som hände mina pojkar . - Till utfrågning . Nu ! Det är en order . 
Kom igen . Hoppa upp . 
Vad glor ni på ? 
Ni har en Flygande fästning att lappa ihop . 
- Fortsätt jobba , pojkar , - Sätt fart ! Kom igen . Sätt fart . 
Starta lastbilen . Inget prat ! Ja . Rena undret att planet inte störtade . 
Nödlandning . 
Motorn var paj . 
Jag måste ta dig till utfrågningen , Buck . Kom . 
Fällde inte en enda bomb . 
Var tvungen att dumpa dem i Kanalen . 
Jag vet . 
Kom nu . 
Varför sa du inget ? 
Vadå ? 
Du har varit uppe . 
Två uppdrag . 
Du berättade inte hur det var . 
Vad skulle jag säga ? 
Du har sett det nu . 
Jag vet inte vad jag såg . 
Trettio killar ... Bara ... 
Jag borde ha varit där uppe med dig . 
Vi har en lång väg framför oss . 
Jag beundrar er amerikaner . Ni bombar i dagsljus . 
Men dagbombning är rena självmordet . 
Du verkar mest vilja strida nattetid , Bryan . 
Vem kan träffa målet nattetid ? 
Känner du inget ? 
För själv känner jag inget alls . 
Vi har problem , major . 
- Jag kan flyga . 
- Så fan heller . 
- Vi leder skvadronen idag . 
Motor tre är illa skadad . Akterskytt till Cleven . Biddick är träffad . 
- Var beredda på kraschlandning . - För lågt . Pilot till besättning . Håll i er . 
