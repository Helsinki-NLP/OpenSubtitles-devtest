Vet att du alltid är i mina tankar , från att jag vaknar tills att jag lägger mig till nattvila . 
Men även då fyller du mina drömmar . 
Du är och förblir den enda flickan för mig . Hoppas jag . 
Uppdraget mot Regensburg-Schweinfurt var vår största och kostsammaste strid dittills med bred marginal . 
Vi miste Biddick , Claytor , Van Noy och deras besättningar . 
Vi visste inte vilka som dödats eller tillfångatagits . 
Där är det tolfte . 
Bättre sent än aldrig , eller hur ? 
Bäst att ha iskall öl redo för pojkarna . 
Räkna inte med det . 
Okej , grabbar , sätt fart . Ja . Hämta er utrustning . 
Vi ska åka hem . 
Nu . 
Mod tog sig många uttryck under kriget . 
För allierade flygare som sergeant William Quinn som hoppade i fallskärm , fanns bara ett sätt att undgå fångenskap . FLANDERN , BELGIEN Hjälp av utländska vänner . 
Den som påkoms med att hjälpa en flygare kastades antingen i koncentrationsläger eller avrättades . 
Riskerna var enorma . 
Sitt här . Jag är strax tillbaka . 
Bailey . 
Du lever . 
Klarade sig nån mer ? 
Ditt är det första bekanta ansikte jag har sett . 
Vem är han ? 
Det är Bob . 
Vilken grupp sa du att du tillhör ? 306:e . 
- Är du skytt ? - Ja . 
Ni måste ha ställt till med ett helsike för tyskarna . 
De gav sig på oss utav bara fan . 
Vi fick vår andel . Nå ? 
Jag har druckit ur en ho sen igår . Och du ? 
Hur gick det med Baby Face ? Och alla andra ? 
Du där . Följ med mig . 
Vad heter du ? 
Sergeant William Quinn . 
Serienummer 6391477 . 
Skriv ner dina svar , tack . 
Vad var ert uppdrag ? 
Att bomba en Messerschmitt-fabrik . Du tjänstgör som ... 
Radiooperatör . 
Skriv ner svaren , tack . 
Gillar du baseball ? Gillar du baseball ? Ja . 
Vilka spelade Babe Ruth för innan Dodgers ? 
Babe Ruth har aldrig spelat för Dodgers . 
Han spelade för Yankees . 
Och före det spelade han för Red Sox . 
Vem står staty på Trafalgar Square ? 
Jag vet inte var det ligger , sir . 
Har du aldrig varit i London ? 
Vi var stationerade i East Anglia . 
Det krävs två dygns permis för att hinna till London . Jag har aldrig haft så lång permis . 
Skriv dagens datum högst upp på pappret . 
Vad heter er nationalsång ? 
Star-Spangled Banner . 
Kan du sjunga den ? 
Jag har inte grillats så hårt sen examen i samhällskunskap . 
Verkligen sant . Jag trodde att jag körde . 
Bob , har du en tändsticka ? Ja . Har du en cigg ? 
Varför sköt du honom ? 
Han var infiltratör . 
Nej , jag pratade med honom i en timme . Quinn ? Du pratade med honom . Han var amerikan . De har försökt infiltrera vårt nätverk på många sätt , men vi avslöjar dem alltid . 
Ni kunde ha tagit fel . 
Vi tar aldrig fel . 
Tjugofem var det magiska antalet . 
Om man överlevde 25 uppdrag blev man hemskickad och fick turnera för krigsobligationer . 
Hur ska pojkarna ta det om Dye inte klarar det ? 
Det blir antingen en sjujäkla fest eller en sjujäkla likvaka . 
På hösten 1943 var kapten Glenn Dye och hans besättning de första som kom nära . 
16 SEPTEMBER 1943 - Pojkar . - Major . Major . Tommy , du kom för att se på . 
Håller killarna dig utanför trubbel ? 
De ställer till trubbel för mig , John . 
Säkert . Billy , Sammy , jobbar ni med de här sluskarna nu ? 
- Såvida du inte har jobb åt mig . 
- Kom och jobba med oss . 
- Gärna . 
- Visst . 
Ena riktiga arbetsmyror , de här . 
Lil , oroa dig inte för Dye . Tjugofem uppdrag . Han är snart här . Tjugofem uppdrag . Han är snart här . 
Tack , John . 
Vi ses , pojkar . 
Hallå där , major . Hallå . 
Du ser ut som en affisch för krigsobligationer . Mycket stilig . Jag känner mig som en sån också . 
- Hej . - Mina herrar . Roligt att höra det från dig , major . 
- Läget , Bucky ? - Jack . Läget ? - Kan inte klaga . - Croz . 
- Major . 
- Hallå . Titta där borta . 
- Det är Dye . 
- Där är han . 
Tjugofemte uppdraget ! 
Du får åka hem ! 
Tjugofem ! 
Du får åka hem , din tursamma jäkel ! 
Han stal din inflygning . 
Han stal din flicka . 
GRATTIS TILL 25 : E UPPDRAGET Vill ni träffa pojkarna ? Följ med mig . 
Där har vi honom . Du verkar roa dig kungligt . 
Akta damen . Akta damen . Nej då . Jag ska ditåt . 
- Hans mamma dog . - Där har vi honom . Vår egen Charlie Robertson . Charlie ? 
Vem är Charlie ? 
1922 . White Sox mot Tigers . Stoppade varenda motspelare hela matchen . 
Siste kastaren som gjorde en felfri match . Tills nu . 
Får du åka hem innan Florida ? Ja . Tre dagar . Kanske jaga med pappa , låta mamma skämma bort mig . 
Sen besöker jag några stationer för att bevisa att det faktiskt är möjligt att klara 25 . 
Ja , med nöd och näppe . 
Det är bara vi kvar , eller hur ? 
Tolv flygbesättningar av ... Trettiofem som flög in från Grönland . 
Det stämmer . 
Vi gläds med dig , Dye . Just det . Vi är glada för din skull . Väldigt glada . Och för killarna som inte är här , men som skulle ha varit det . Och för killarna som inte är här , men som skulle ha varit det . 
- Skål för dem . - Ja . 
Ja , skål för dem . 
Mina herrar , jag ska se till pojkarna , så att de inte firar för hårt utan mig . 
- Charlie Robertson . - Vad försöker han göra ? 
En klar . 
Sluta stirra . 
- Jag stirrar inte . 
Gjorde du ? Nej . Är ni inte bekymrade alls ? 
Jo , jag är verkligen bekymrad . 
- Det är Nash . Han är som han är . - Nej , jag menar inte det . 
Jag menar att vi har en jättefest för att en av oss inte åker hem i likkista . 
Varför ? Varför säger du jämt såna saker ? 
Titta vem vi har här . 
Se upp , killar . Här kommer danskungen . 
Nej , uppmuntra honom inte . Han skrämmer bort damerna . 
Fin stil . 
Mina herrar , vad har jag missat ? 
Jag spanar in brudar , och Farsan här försöker sänka stämningen . 
- Med andra ord , ingenting . - Dämpa . Stämningen . Du menar " dämpa " stämningen . Stämningen . Nej . Jag sa bara att det är ett dåligt tecken för oss . 
En besättning överlever , och man har en jättefest ? 
Alla piloter gör så . - Du vet att de är på dig , va ? - Det hoppas jag . 
- Killar ? 
- Mina herrar . - Major Egan . 
Major Cleven . 
Rosenthal . Nash . 
Det stämmer . 
Andrepiloterna , Spatz and Lewis ? 
- Speas . Sir . - Speas . 
Lewis , sir . Men alla säger Farsan . 
- Okej . - Hör ni , killar ... Var ni piloter före kriget ? 
- Jurist , sir . - Jurist ? 
- Var lärde du dig flyga ett B-17 ? 
- Laredo . Nio månader , 12 timmar dagligen . - Mm . 
Skytteutbildning . Löjtnant Nash också . 
Tja , pojkar , ert rykte föregår er , ska ni veta . 
Menar du att vi flög i undertröjorna , sir ? 
Jag hänger inte med . 
Vi var kända för att flyga i underkläderna . 
Ni allihop ? 
Ja , sir . Är det så ungdomarna gör nuförtiden ? 
I Texas blir det så hett i planen att man kan steka ägg på instrumentpanelen . 
Verkligen ? 
Vi hade inte hört om underkläderna , men vi hörde att ni är utomordentliga piloter . 
Vi är glada att tjänstgöra i kriget , sir . 
Vi har ansökt om stridande position i flera månader . 
Nu när vi är här , känns det som om vi faktiskt ska uträtta nåt . 
Nog ska ni uträtta nåt , allt . 
- Roa er nu . 
- Ja , sir . 
- Gosse . Varför måste han nämna det där ? 
- Vad tänkte jag på , som pratar om mina underkläder inför ... 
- Ingen fara . - Be för mig . Jag tar chansen . 
Löjtnant Herbert Nash . 
Helen . Som Helena av Troja . 
Inte reste du väl runt halva jordklotet för att dela ut kaffe och munkar ? för att dela ut kaffe och munkar ? 
Jag ville göra en insats , och så här blev det . 
Otur för dig , med de här . Jag klagar inte . 
Du ger väl såna blickar till varenda basse som vill ha frukost . 
Nåja ... jag kanske är det sista söta ansikte de nånsin ser . 
Men hur ska jag kunna veta ? Veta vadå ? 
Om du tycker synd om mig eller om du vill kyssa mig . 
- Du gillar nog hennes leende , Buck . - Major Egan . Major Cleven . 
Jag hörde att ni redan har flugit tjugo uppdrag . 
På ett ungefär . 
Han har flugit tjugoen . 
Några goda råd ? 
Försök hålla dig vid liv . 
Under minst elva uppdrag . 
Jaha . Vad händer efter det ? Då har du överlevt det värsta . Eller också inte . Du förstår ? 
Tack , major . Major . - God natt med dig . 
- Tack detsamma . 
Alla de här är nya ansikten ... Om vi störtar blir vi inte heller hågkomna . Som om vi inte funnits , Buck . 
Spelar det nån roll ? Nej , antar jag . 
Mina killar . Överste Harding . Lyssna . 
Jag hade just ett trist samtal med Doc Stover . 
Han tror att ni mjukisar kan bli skjutglada . Han tror att ni mjukisar kan bli skjutglada . 
Inte vi inte , sir . 
Jag sa åt honom att det här är krig och ju längre man är i elden , desto mer tär det på en . 
Så har det varit ända sen den första jädra grottmannen tog en klubba och gav sig på en annan . 
Gick grottmän i terapi ? - Nej . - Inte vad jag vet , sir . 
Verkligen inte . 
Det som räknas är att ni är redo för strid när det gäller , visst ? 
Vad ni gör däremellan ... - Jag gillar er stil , sir . - Jajamän . 
Sån här luftkrigföring fanns inte på grottmännens tid , sir . 
Givetvis inte , Red . Varje krig innebär förändringar . 
Vem tusan gjorde dekorationerna ? 
Jag satte ihop en kommitté , sir . 
Det jädra planet verkar vara på väg att störta . 
Avskeda kommittén . 
Nästa gång bryr jag mig inte . 
Kom , samlas här . Jag har nåt att säga till er . Kom , samlas här . Jag har nåt att säga till er . 
Vet ni hur vi kan göra slut på kriget redan ikväll ? Vi fyller en Flygande fästning med så många bomber som ryms , och pulvriserar Hitlers jävla gömställe . 
Red och Bubbles kan säkert lokalisera den mustaschprydda lilla fan . 
Ja , sir . 
Vem är det nu som är skjutglad ? 
Vem ? 
Ni . 
Nej , du . 
Nej , ni . Sir . 
Lediga ungston . 
Kom igen , pojkar . Nu går vi till aktion . - Lediga ungston . - Order är order . - Sätt igång , mannar . - Hallå , Tatty . 
Du kan inte stå emot . - Gratulerar . - Du kan inte stå emot . 
Du behöver ledighet . 
Översten borde ordna en helgpermis åt dig . 
Du borde följa med . 
London . Kom igen , Buck . Vi gör stan . 
Jaha , kanske nästa gång . 
Hit , Meatball . 
Vill du dansa ? 
Jag skvallrar för Marge , Buck . 
När jag gick ut i kriget var det sista jag väntade mig att tillbringa en månad på en belgisk bondgård . att tillbringa en månad på en belgisk bondgård . 
Vi har fler nedskjutna flygare än tillförlitliga guider . 
Jag vet . Jag tillhör de tursamma . 
Men inte som han . Kom nu ! 
Kom , Romeo . 
Hej , broder . 
Vart tror du att de tar oss ? Nån aning ? 
Vet inte . Via Frankrike in i Spanien , antar jag . 
Ja , jag undrar . Och om vi nånsin får träffa kamraterna igen . 
Alice dök ganska tvärt , så jag tvivlar på det . 
Men Hinton hoppade . 
Ja , absolut . Baby Face hittade nog en utväg . 
Tyst . 
Är hon din dotter ? 
Michou är er guide . 
Hon är bara barnet . 
Hon är er guide , och ni ska göra som hon säger . 
Vad sa hon ? 
Jag vet inte . 
Ge mig den nu . Vadå ? 
Lägg av . Det där behövs inte . 
Om tyskarna hittar den här , vad tror ni att de gör med Louise och hennes familj ? 
De torterar dem tills de talar . Och när de har namnen de behöver , skjuter de dem . 
Sen hittar de nästa och gör likadant med dem . 
Som att repa maskor av en tröja . 
Jag ... Förlåt mig . 
Det var dumt av mig . 
Vad betyder det där ? 
Här betyder dumhet döden . 
Så , hur hamnade du i London ? 
Med drinken köper du småprat , inte en sorglig levnadssaga . 
Jag visste inte att jag köpte nånting alls . 
Tänker du inte försöka få mig i säng ? Tänker du inte försöka få mig i säng ? 
Jag har inte tänkt så långt än . 
- Jag antar att om du ville köpa ... - Mm . ... kunde du hitta nån i Piccadilly . 
Du behöver inte komma ända till Hammersmith . 
Är det där jag är ? 
Major i flygvapnet , men ingen navigatör . 
Nej , pilot . 
Gissa hur man vet om nån är pilot ? 
Hur då ? 
Han lär berätta det . 
Min man är pilot . 
Så du är gift ? 
- Hur länge har du varit soldat ? 
- Sen före kriget . 
- När lämnade du Polen ? 
- När tyskarna invaderade . 
Ja , jag såg journalfilmerna . 
Det var därför jag tog värvning . Före Pearl Harbor . 
En amerikansk hjälte . 
Jag kanske var ute efter äventyr . 
Var är maken ? 
En del piloter överlever för att strida igen . Han stannade kvar . 
Han ville bli hjälte , som du . 
I fjol träffade jag nån från hans skvadron . 
Han sa att Pavel sköts ner över Schlesien första veckan . 
Han är antingen krigsfånge eller ruttnar i en potatisåker . 
Kanske kommer den här spriten därifrån . 
Vill du hoppa i säng med mig ? 
Låt oss dansa först . 
Jag har aldrig varit på mottagarsidan av en bombning förut . 
Mottagarsidan . Märkligt ord för döden . 
Jag har fällt många bomber . Troligen dödat många människor . 
Vilket jävla jobb . 
Känner du dåligt samvete ? 
Gör inte det . Tyskarna förtjänar varenda en av era bomber . 
En del anser att det är skillnad mellan krig och vettlöst mördande . 
Men inte de . 
Vad anser du ? 
Att vi ska vara lika skoningslösa och hårda som de var mot mitt folk . 
Det vore rättvisa . 
Ja , men om det handlar om balans , är mitt öde beseglat för länge sen . 
Det finns ingen balans . 
En händelse följer på en annan . 
De sämsta klarar sig oskadda . De sämsta klarar sig oskadda . De oskyldiga dör . 
Men vet du en sak ? Ju närmare döden man är , desto mer levande känner man sig . 
Varje sekund är en smula död . 
Och jag som tyckte att jag blir teatralisk när jag dricker . 
Vi ses där uppe , Buck . 
- Vi bockar av ett uppdrag till . - Ja . 
Lycka till , kompis . 
Vill du ha en munk ? Nej . 
- Tack . - Den är varm . Försiktigt . 
- Kaffe till , löjtnant ? 
- Har du saknat mig ? 
- De fyra timmarna sen vi sågs ? 
Nåja , det här blir längre . 
Hur ska jag stå ut ? 
Vad är det ? 
Du kanske är den sista söta flicka jag nånsin ser . 
Säg inte så . 
Och du är ta mig tusan den sötaste . 
Vi ses senare . 
Absolut . 
- Titta , vår egen Adonis . - Lägg av . 
Vårt första försök att bomba Bremen var en katastrof . 
Men det kändes som en livstid sen . Vi var redo att försöka bomba de där ubåtsbaserna igen . 
Ingen var mer redo än major Cleven . 
Funkar den ? 
Nej . Jäklar . 
Major , jag har problem med vänster magnetspole i motor två . Den ger ojämna pulser . 
Det är nog bara brytarspetsarna . Jag fixar dem medan ni startar . Tre motorer ? 
Jag klarar det , sir . 
Galet . Tänker du följa med runt ? 
Gör ett försök . 
Jag vet inte , Buck . 
Att laga en magnetspole på startbanan är en sak . Men i rörelse ? 
Om Lemmons lovar att fixa det , så gör han det . 
Du måste ha tro . 
Hur går det , Lemmons ? 
Vi måste leda skvadronen . 
Jag håller på , major . Jag jobbar så fort jag kan . 
Vi har två plan kvar , Buck . 
Vi har två plan framför oss . 
Ja , sir . 
Ett plan kvar , Buck . Det är nu eller aldrig . 
- Ett plan kvar , Lemmons . 
- Det är inte för sent att avbryta , Buck . - Vi kan köra till höger där borta . - Vi leder skvadronen . 
- Vi leder skvadronen . 
Kom igen , Lemmons . Sätt fart . 
Nu kan ni flyga . 
Nu kör vi , pojkar ! 
DeMarco , erkänn att du hade fel . Okej , jag hade fel . Nu kör vi . Okej , jag hade fel . Nu kör vi . Jajamän , kör ! 
PARIS , FRANKRIKE På stationen finns det många tyskar . 
Gör som jag gör . Om jag tar fram mina ID-handlingar gör ni det också . Om jag tittar på klockan gör ni det också . 
Vad ni än gör , tala inte . 
Förstått ? 
Ska vi gå ? 
Nej , jag ska gå på toan . 
Nu ? 
Tror du att de skiljer oss åt ? 
Jag vet inte , Bailey . 
Jag måste fråga dig en sak , Quinn . 
Det har gnagt på mig . 
Beträffande kraschen . 
- Är Baby Face ... 
Jag fick inte loss honom . 
Spaken satt fast . 
Jag försökte verkligen . 
Jag lämnade honom kvar . 
Lilla Baby Face . 
Jag försökte . 
Jag vet inte . 
Jag hade också hoppat . 
Biljetterna , tack . 
Och ha era papper klara för myndigheterna på stationen . 
Nej , herrn , det är för myndigheterna . 
Era biljetter , tack . 
Ett ögonblick , herrn . 
Ursäkta mig . - God dag . - God dag , fröken . Biljetten , tack . 
- Här . - Här . 
- Tack . 
Biljetten , herrn ! 
Herrn , jag behöver se er biljett ! 
De är döva . De hör er inte . 
Titta i era fickor ! 
Vad är det med er ? De är döva . Han förstår inte . - Varför flyr han ? 
- Han blev rädd . Tänk er själv . 
Vänta . 
Stanna . 
Du måste vända dig om och gå lugnt tillbaka till kupén . Förstått ? 
Har ni er biljett ? Ja . 
Ta fram den . 
Har ni hittat biljetten ? - Konduktören ? - Ja , fröken ? Nån har stulit väskan för en stackars dam ! 
Ja . Ett ögonblick , fröken . 
Sätt er och behåll lugnet . 
Tänker ni inte göra nåt ? Tänker ni inte göra nåt ? Lugn . Nåväl . 
Där borta . En liten tjuv ! Titta . Han är rödhårig . 
Gör inte om det där . Förstått ? 
Har du varit här hela tiden ? 
Det här är Manon . 
Vi har en lång väg kvar . 
Vi ska ta er till Spanien och hem till England . 
Men ni måste behålla lugnet . 
Om du gör om det där , knockar jag dig . 
Dra inte till för hårt . 
Lämna startbanan . Jösses . Sätt fart ! Var redo , pojkar . Lämna startbanan . 
Elva , tolv . - Tretton . - Tretton . 
De är tretton . 
Var är du , Buck ? 
- Inga fler . - Ja , sir . 
Vi hade tjugofyra bombplan . Tretton kom tillbaka . 
Tre med motorfel . Sammanlagt åtta som vi miste . 
Det blir åttio man . 
- Sir . - Några ersättare . 
Kidd och Blakely . 
DeMarco och Buck Cleven också . 
Sir . Löjtnant Crosby ? 
Jag beklagar . 
Förbannelse över Bremen . Buck . 
Vad är det ? 
De klarade sig inte . 
Vem ska ta hand om Meatball ? 
Låt mig hjälpa till , doktorn . 
Rosie ' s Riveters . 418:e . 
- Varsågod . - Tack . - Allt väl ? - Skönt att ha er tillbaka . 
- Här finns kaffe . - Kaffe på den sidan . 
Kom . 
Det var som att flyga genom en solid mur av luftvärnseld . 
- Fortsätt . - Ett FW körde rätt in i dem . - Fortsätt . - Ett FW körde rätt in i dem . Båda planen sprängdes . Hur var förhållandena ? Kunde ni se målet ? 
- Skvadronledaren störtade . Hoppade nån ? Såg du några fallskärmar ? 
Jag såg fyra fallskärmar . Inga fler . 
Jag förstår . Hur skildes ni från gruppen ? 
Det var så förvirrat där uppe efter att ledarplanet för 350:e störtade . 
Vårt plan med Buck Cleven och DeMarco . 
Hela första avdelningen . 
Nash och Speas också . 
Jag såg inga fallskärmar . 
Vänta lite , Farsan . 
Helen . 
Det var ett helvete där uppe idag . 
Löjtnant Nash överlevde inte . 
Jag beklagar . 
- Crank . - Hallå . Såg du hur det gick med Blakelys och Croz plan ? När ? Var ? Hur många fallskärmar ? Nej , de lämnade formationen nånstans vid referenspunkten . 
Och Buck ? 
Vem berättar för Egan ? 
God morgon . 
Morgon ? Klockan är över tolv . 
Återställare . 
Jag har huvudvärk . 
Nej , du behöver en återställare . 
Det är boten . Jag måste gå . 
Har du bråttom nånstans ? 
Vi ska inte göra mer av det här än vad det var . 
Det var jäkligt bra . Hur kan det bli bättre ? 
Du , jag ska gå ut idag och få nåt att dricka . 
Jag ska roa mig . Jag skulle gärna göra det med dig . 
Mitt hjärta klarar inte ännu en död pilot . 
Jag vet att du förstår raring . 
Ursäkta , vet ni var man kan köpa en dagstidning ? 
Där borta . Runt hörnet . 
Herregud . 
Låt mig se henne . Gode Gud . - Tack . 
Låt mig se henne ! Är hon död ? Nej , det är hon inte ! 
- Behåll växeln . 
Norfolk 7322 , tack . 
- Bowman här . 
- Red , Egan här . 
Hur gick matchen igår ? 
Inte så bra som vi hoppades . 
Var Buck med i matchen ? Ja . 
Spelade han bra ? 
Han gav allt in i det sista , John . 
Vilka fler ? 
De flesta i förstauppställningen . 
Blir det match imorgon ? Ja . 
Okej , hälsa coachen att jag ska vara där i tid . 
Och , Red jag vill leda laget . 
I NÄSTA AVSNITT Ni behöver inte undra . 
Ni förstår allihop varför jag kom tillbaka i förtid . 
Ett nytt uppdrag . 
Målet är strax öster om stadens centrum . 
Det är mycket folk i katedralen . 
Vi har aldrig bombat så nära - civila befolkningscentra förut . - Jösses , Crank . Det är krig . Vårt jobb är att fälla bomber . 
Jag fick den igår . Men den flyger nog . Då är jag helt lugn . 
Jaktplan klockan tolv . Jösses . 
Motor ett stannar . 
Motor fyra stannar ! Motor fyra stannar ! 
Vi måste komma härifrån fort . 
Vet du när min bombgrupp landar ? 
Var är våra pojkar , Chick ? 
