Länkar till S-band 4 . 
Signalen är låst . 
Okej . Vi är inne igen . 
Redo att sända krypterat testping till Ranger . 
Kolla att han fick rätt kryptering . 
Måtte det funka nu . 
Jag tror på det här . 
Det har du sagt 20 gånger nu . 
Nitton . 
Sändtagare uppkopplad . 
Kringgår säkringen . Ping . 
Sänder ping till Ranger . 
VERIFIERING NEKAD Nix . Deras detektor nobbade oss igen . 
Sam har varit ombord på Ranger i en månad . Hon borde ha satt dit vår vid det här laget . 
Om hon inte kopplar in vår detektor inom 48 timmar ... Så går Guldlock mot jorden . Och det kan vi inte göra nånting åt . 
Ranger , Happy Valley . Sänder simulerad order om motorstopp . MOTTAR Bekräfta mottagande och autentisering . 
Happy Valley , Ranger har just mottagit er simulerade order om motorstopp . 
Huvudmotoravstängning verifierad vid 19 minuter och 58 sekunder . 
Och motorn signalerar avstängning . 
Snyggt gjort , Ranger . Det var tjusigt . 
Det behövs bara överlägsen slughet och skicklighet , kommendör . 
Vi kör övningen igen om sju timmar . 
Vi måste få in drillen . Vi får inte en andra chans i skarpt läge . 
Uppfattat , Happy Valley . Vi kör igen om sju timmar . Klart slut . 
Klart slut . 
Okej , gott folk . Vi fortsätter med nedstängningssimuleringen . 
Verifierad detektor aktiv ? 
Detektorn signalerar aktiv . 
Ställ ner uteffekt till reservläge för fusionsreaktorer 1 till 4 . 
Fusionsreaktorer 1 till 4 i reservläge . 
Bra . 
Rozhenkova , simulera 50 % termaleffektreduktion på reaktorer 1 till 4 . 
Simulerar 50 % effektreduktion på reaktorer 1 till 4 . 
Mr James , vänligen rapportera om vår mekaniska infästning i asteroiden . 
Ankarpåfrestning nominell på alla punkter . 
Sensorisk självkontroll visar inga fel . Allt klart . 
Utmärkt . 
Framdrivningssystemen nominella . Temperaturer och tryck inom toleransen . 
Okej . Vi kör en simulation med för högt tryck på argontank 2 . 
Primära och sekundära . 
Bekräftar . 
Jösses . Den är rökt . Inga kontrollsignaler från NASA kan passera genom den här . 
Vi har inte tid att laga den . Nästa borrning är om tre timmar . 
Logga felet . Sätt in reserven . 
Jag vet var den finns . Jag hämtar den . 
Tack , Massey . 
Detta är metankoncentrationerna robotarna upptäckte vid testet i lavatunnlarna precis utanför Happy Valley . Och detta är data de skickade i morse från Korolevkratern . 
Det är förstås bara preliminära resultat , men ... Dev . 
Förlåt . 
Är det där Korolevkratern ? 
De största koncentrationerna finns där , ja . Men det kommer också tydliga signaturer från Chasma Australe nära sydpolen . Ingendera regionen är känd för vulkanisk aktivitet . 
Några data än om vad som producerar metan ? 
Möjligen vulkanisk aktivitet djupt under ytan . Eller ännu bättre , högsta vinsten . 
Metanogena bakterier ? Liv . 
Då har du lite att stå i . 
Okej . Fortsätt , Kelly . Om det finns liv på Mars , vill jag att du är den som finner det . 
Ska du gå ? 
Jag har mycket mer data att visa dig . 
Jag är strax tillbaka . Jag måste ordna några saker . 
Med min pappa ? 
Varför frågar du ? 
Ni har tillbringat mycket tid tillsammans på sistone . 
Vilket faktiskt är förvånande med tanke på er historia . 
Ja , han ... Hans erfarenhet här uppe är otroligt värdefull inför infångningen av asteroiden . 
Han nämnde inte att han jobbar på det . 
Men jag har ju inte sett honom på några dagar , så ... Ja , det har varit mycket tidskrävande . Men han är glad att ha er här . Han pratar jämt om den där lilla pojken . 
Ja , jag ... Bra att de finner varandra . 
Jag trodde bara ... Jag vet inte . 
Att även vi skulle vara närmare . 
Det låter väl dumt med tanke på allt som ... Inte alls . 
Jag förstår . Tro mig . 
Jag fick aldrig chansen att försonas med min pappa . 
Men du har ännu chansen . 
Jag måste gå . 
Du . Bra jobbat , Kelly . 
Vill ni ha våra övervakningskameror ? 
Vi måste se hela basen , så att ingen kommer på vad vi gör . 
Farligt . Det är mycket farligt . 
Liksom att vara ensam i en nordkoreansk kapsel i sju månader . 
Det var inte ett val . Men detta är ett val . 
Min fru . 
Vad är statusen ? 
Lee , det är komplicerat . Berätta . Hon är i fara . 
Som jag sa förut rör det på sig . 
Vi har en bra plan för att få henne ut ur Nordkorea , men att smyga henne ombord på en Heliostransport är ännu mer komplicerat . 
Lee , inser du inte vad vi gör här ? 
Den här asteroiden kommer att säkra framtiden för Mars , för dig och din fru . 
Det är bra att ha sin familj hos sig . Som du har . 
Jag ska hjälpa . 
Bra att ha dig med ... Okej . Jag får video och ljud från PRK . 
Och nu har vi Op-centralen . 
Jag trodde aldrig att jag skulle säga det här , men Gud välsigne Nordkorea . 
Redo för statusuppdatering ? 
Reda att länka när ni vill . 
Happy Valley , bekräftar att vi har reservdetektorn installerad i god tid före nästa simulering . 
Hörde ni ? 
Samantha Massey verkar ha levt upp till mina förväntningar . 
Uppfattat , Ranger . Tack för uppdateringen . 
Men för säkerhets skull testar jag igen . 
EECOM , förbered nästa simulering för överföring till Ranger . 
Skicka ett ping till . 
- Vi är inne . - Ja . - Kom igen . Ja . - Ranger godkände vårt ping . 
Bra jobbat , allihop . 
Vår detektor är installerad och vi styr maskinerna . 
Då kör vi . 
Och efter många riskbedömningar den senaste månaden , kan vi inte utvidga brytningsschemat mer . BUDGET OCH TIDSSCHEMA Presidenten kommer att bli besviken över att det tar två år tills vi har en färdig produkt . 
Det måste finnas ett sätt att få fram säljbart iridium fortare . 
Vi kan bygga fler skepp , borrar , lastmaskiner . 
Det kommer dock att driva upp kostnaderna . 
Jösses , nej . Vi talar redan om en triljon dollar . 
Om jag säger åt honom att det blir ännu dyrare , kanske han avskedar oss alla . 
Nåja , tack för era tankar . 
Fortsätt kläcka idéer , så kanske vi hittar nåt som funkar . 
Okej . Eli , när kan vi vänta oss grönt ljus för anslag till nästa generation Marsfarkoster ? 
Låt mig återkomma om det . 
Men vi närmar oss vår tidsgräns . 
Tänk bara vad vi skulle kunna åstadkomma om inte de där jävla politikerna var i vägen . 
Det enda de är bra på är att uppskjuta beslut tills absolut nödvändigt . 
Kan jag få din åsikt om de här kalkylerna för projektilbanan ? 
Ge det här till Sergei . 
Jag vill att nån mer tittar på de här projektilbanorna . 
Vi måste vara helt säkra på att vi har räknat med värsta tänkbara scenario innan vi går till dem som bestämmer . 
Nej , det får vara nog . 
Jag har förmedlat anteckningar mellan er den sista månaden . 
Vi har inte tid med denna snigelkorrespondens . 
Men vi behöver hans hjälp . 
Han förstår projektilbanor bortom månen bättre än nån annan . 
Okej . Men det måste ske ansikte mot ansikte . 
Var ? 
De bevakar mig dygnet runt . 
Vi kan mötas hemma hos mig . 
Vi säger att vi jobbar på det här . 
Det är riskabelt . 
Säg nåt som inte är det . 
- Det är fel på bildskärmen . - Va ? 
Den har inte varit statisk förut . 
Det kanske är en gammal monitor . 
Vad pågår ? 
Övervakningsmonitorerna fallerar . 
Klart att de fallerar . Rena eländet ! 
Sir , låt oss lösa problemet , ni ska inte behöva ... Vänta lite ... 
Vad är det här ? 
Jag vet inte . 
Denna amerikanska spionutrustning hittades på Demokratiska folkrepubliken Koreas territorium ! 
Vi kräver en förklaring till denna skandal ! 
Så ni fann den här i ert komplex ? 
Den gör bildskärmen statisk . 
Vilken bildskärm ? 
Hon frågar vilken bildskärm . 
Jag förstår . Den var inkopplad på systemet ni använder för att spionera på oss . 
Säg att den Demokratiska folkrepubliken kräver att den skyldiga ska straffas ! 
Befälhavare Cho kräver att ni utreder . 
Jag hjälper gärna till , men i så fall måste vi få tillträde till ert komplex för att se var apparaten upptäcktes . 
Hon vill att hennes folk får genomsöka vår modul . 
Nej ! 
Ett intrång på Folkrepublikens område kommer att få svåra konsekvenser . 
Jag har inte tid med det här just nu . 
Kan det vänta tills efter asteroiduppdraget ? 
Kommendören ber om ursäkt för olägenheten . 
Under tiden kan jag spåra dess ursprung . Den har ett NASA-serienummer . Mer kan jag inte göra just nu . 
Hon ska vidarebefordra era krav till NASA . 
Hon förhalar . 
Säg åt henne att genast gripa och förhöra Helios tekniker Miles Dale . Bara han har varit i vår modul . 
- Befälhavaren vill uttrycka sitt ... - Miles Dale ? 
- Ms Talmadge ? - Ja , kommendör . 
Jag vill att du spårar en apparat . Varifrån den kom , vem som hade tillgång . Genast . 
Ska bli . 
Hon är ett värdelöst redskap för det dekadenta kapitalistsystemet . 
Jag ska undersöka saken själv . 
- Tack . - Du , Lee . Hur mår du annars ? 
Hur mår Moon Yeong ? 
Det är jobbigt att vara isär . 
Ja , jag vet vad du menar . 
Men vi är snart tillbaka på jorden . 
Vet du , Zay , av allt jag har gjort i livet är jag mest stolt över dig . 
Att se dig växa upp och bli en fin ung man som nu har en egen familj . Jag bara ... Det betyder mer för mig än nån utmärkelse i världen . 
Och jag tänker bli världens bästa farmor . 
Så , tre månader till den stora dagen , va ? 
Ja . Då borde Guldlock vara på väg mot jorden . 
Liksom jag . 
En sak jag sörjer över är att jag inte fick se dig ta dina första steg eller säga dina första ord . 
Men nu får jag se din dotter göra det . 
Förlåt , det ... Det tog mig med överraskning . 
Jag är bara så lycklig . 
I alla fall ... Jag vet att du avskyr Star Trek , men bäst att du vänjer dig , för jag tänker se till att mitt barnbarn blir en fanatisk Trekkie . Just det . Vi ska se alla säsongerna . Alla tre . 
Och Twilight Zone , och Bob Newhart Show . 
MASH , Columbo ... Margo . 
Kom in . 
Tack . 
Är ... Jag kom hit för några timmar sen . 
Och ingen såg dig gå in ? 
Jag parkerade långt bort , gick över grannars tomter . 
- Tack för att du kom . - Självklart . 
Ska vi börja ? 
Med dessa uppdaterade CG-uppskattningar kan vi beräkna drivkraftvektorerna . 
Man behöver också beräkna masscentrumspridningen . Från tröga kompressionskrafter under starten . 
- Väldigt smart . - Instämmer . 
Med projektilbanan inställd kan vi börja gruvdrift på Guldlock inom nio månader . 
Det är positivt , ja . Men det är ändå synd . 
Vad menar du ? 
Asteroiden kommer till jorden och alla investeringar med den . 
Det finns inte längre skäl att satsa mer pengar på Mars . 
M-7 har ett starkt åtagande på Mars . 
- De sa ... - Ja , det de alltid säger . 
Men Korzhenko bryr sig bara om att berika sig och sina kumpaner . 
Nu kommer asteroiden att göra det , och de kommer att lämna Mars åt sitt öde , och NASA gör likadant . 
Precis som de gjorde med Marsprogrammet på 80-talet . 
Tills vi gjorde det nödvändigt . Minns du , Margo ? 
Utan konkurrens , inga framsteg . 
Det får räcka med geopolitiskt skoj för i kväll . 
Barn , ta bort tallrikarna . 
- Förlåt att vi kapade ditt hem , Victor . - Ingen fara . Det är okej . Fortsätt ni . Barnen måste i säng . 
Pappa , klockan är bara nio . Jag vet . Kom nu . 
Innan du går , här är nånting gott . 
Tack . 
Tack . 
Margo . Jag har en sak till dig också . - Glöm inte att borsta tänderna . - Jag har inte hört den skivan sen alltför länge . 
Har du ... Har du tänkt mer på min idé ? 
Att vi sticker ? 
Jag ... Jag har inte hunnit . 
Vi har så mycket kvar att göra . 
När asteroiden väl har kurs mot jorden kommer Irina Morozova att beordra dig tillbaka till Moskva , 
Det ... Det vet du inte . Det kan bli fler tillfällen . 
Nej , det kan det inte . 
Så vad gör vi ? 
Vi sticker iväg , gömmer oss i en lägenhet nånstans och glor på väggarna de kommande 20 åren ? 
Jag har en högt uppsatt vän i det brasilianska rymdprogrammet . 
Vi tar kontakt med honom och erbjuder våra tjänster i utbyte mot regeringens beskydd . 
Skulle de gå med på det ? 
De skulle vara överlyckliga . 
Du och jag kan göra Brasilien till en stormakt i rymden . 
Som den första tiden med Apollo-Soyuz . 
Jag föreslår Soyuz-Apollo , för enkelhetens skull . 
Tillsammans ska vi fullborda det vi påbörjade . 
Jag måste tänka på saken . 
Vi har så lite tid , Margo . 
Jag vet . Men jag måste få det här uppdraget i hamn först . 
Videoserienumret som ni kan se här , visar att komponenten anlände till Phoenix med den senaste transporten . 
Den registrerades här . Det finns inga uppgifter om att den lämnat Phoenix . 
Och den lastansvariga fann kartongen där den skulle vara enligt inventarielistan . 
Sigillet var inte brutet , men när hon öppnade kartongen hade innehållet bytts ut . 
Eli , du håller säkert med om att detta visar på ett allvarligt problem . 
Senaste inventeringen var för en månad sen . 
Personalen skannade bara förpackningarna . De kollade inte att innehållet matchade etiketterna . 
Jag beordrade en noggrann inventering , som avslöjade många stölder främst kommunikations - och datorutrustning som du ser i den bifogade filen . 
Eli , vi har nog att stort problem här . 
Inte bara stölder , utan kanske nåt mycket allvarligare . 
Jag menar , vad ska de använda den där utrustningen till ? 
Skicka hit Will Tyler . Och be Irina Morozova i Moskva att kontakta mig . 
Befälhavare Cho , ert te är klart . 
CIA har granskat listan med stulen utrustning . 
Det är avancerad kommunikationsutrustning utan värde på svarta börsen . 
Så varför stjäla den ? 
Enda syftet är att övervaka och kommunicera med en rymdfarkost . 
Den enda rymdfarkosten som fraktar last med avsevärt värde - i Mars närhet är ... - Ranger . Helvete ! 
Med tanke på sabotagen i Happy Valley nyligen måste vi se mycket allvarligt på detta hot . 
Tror du att nån vill sabotera asteroiduppdraget ? 
Vi måste anta det . För mycket står på spel för att blunda för det . 
Här är vi nu , redo att förvandla liven för sex miljarder människor till det bättre och en handfull anarkister vill förstöra alltihop . 
- Varför ? 
- Som Dostojevskij sa en gång : Om man bygger att palats av kristall , oavsett hur vackert , finns det alltid någon idiot som vill rasera det . 
Det är förstås lite förenklat . 
Nåja , vilka det än är måste vi hitta dem innan de utför sabotage mot Ranger . 
Vi har bra folk ombord på det skeppet , och inga fler liv får gå förlorade så länge jag bestämmer . 
Det är mindre än 24 timmar till start . 
Om de tänker göra nåt , agerar de innan dess . 
Jag rekommenderar att aktivera våra hemliga agenter i Happy Valley för att samla mer information . 
Låt CIA och KGB ta reda på vilka som ligger bakom . 
Tim , ring upp direktor Hanlin . 
Inte förvånande att det finns underrättelsepersonal här uppe , men Mike , jag trodde aldrig att du var en av dem . 
Om du gjorde det , vore jag usel på mitt jobb . 
Och mr Avilov . Alltså , du var rätt aktiv under strejken . 
En agent måste smälta in i mängden som fiskarna i havet . 
Så , jobbar KGB och CIA hand i hand nu ? 
Precis som ni gjorde på Apollo-Soyuz . 
Ja , det var mycket modigt . 
Vi vet alla hur viktig Guldlock är för våra två länder . 
Därför måste vi gå till botten med det här . 
Folks liv står på spel . Folk vi alla känner uppe på Ranger . 
Vi har några idéer om var vi ska börja . Bra . En sak till . 
Nordkoreanerna nämnde nån Miles Dale för mig . Det kanske är ett blindspår . 
Jag känner till honom väl . 
Han säljer på svarta marknaden . 
Han kan vara inblandad . 
Bra att veta . Vi ska prata med honom . Bra . Håll mig underrättad . 
Under tiden godkänner jag ännu en genomsökning av basen . 
Pappa ? 
Kel . 
Hej , pappa . 
Hej . Är allt okej ? 
Vi måste prata . 
Jag är ledsen , raring . Jag ... Jag kan inte nu . Så ... - Varför inte ? 
- Jag kan bara inte . Det är en sak med jobbet , så ... Ja . 
Ja , jag vet . Team genomsöker hela basen efter saknad kommunikationsutrustning . 
- Ja . - Vet du nåt om det ? 
Nej . Varför skulle jag det ? 
Jag vet inte . Du tyckte förut att Dev Ayesa var ondskan i människohamn . 
Nu är ni plötsligt bästa kompisar och viskar i hörnen . 
Kan du inte berätta vad som pågår ? 
- Inget pågår . Jag lovar . - Sluta ljuga för mig . 
Du tror att jag inte märker nåt , men jag känner dig , pappa . 
Du har ljugit för mig ända sen jag kom hit . 
Innan dess också . 
Vad är det egentligen med dig ? 
- Vart ska du ? - SL3-14 . Systemreparation . 
Fortsätt . 
Kom in . 
Hejsan . Jag är här för att laga luftcirkulationen . 
Skönt att höra . 
Ja , vi har ett stort problem . 
Men inte med luftcirkulationen . 
Sätt dig . 
Som ung var jag inte rädd för nånting . Inte ens döden . 
Jag trodde alltid att jag skulle dö som en hjälte . 
Gordo . Han berättade en gång om sin pappa som fick cancer . 
Pappan var marinsoldat . Tuff som tusan , men mot slutet var han skräckslagen . 
Jag bara ... Jag vill inte sluta så , Kel . 
Skälet till att inte komma hem var att jag inte vill sluta på ett vårdhem med blöja och dregelskydd , klämmande på en boll framför tv:n och inte minnas vem fan jag är längre . 
Här uppe gör jag nåt meningsfullt . 
Jag bygger nånting . Nåt som kan vara långt efter att jag är död . 
Kanske hans barn också . 
Varför berättade du inte det här förut ? 
Du skulle väl tro att jag var knäpp . 
Jag tror inte att du är knäpp . 
Kanske bara lite . 
Jag är ledsen , Kel . 
Jag borde ha funnits där för dig och Alex . 
Och jag borde inte ha ljugit för dig . 
Aldrig . 
Så tänker du berätta vad du och Dev har i görningen ? 
Radioapparater , kablar , nätverkskopplingar , monitorer . 
Flera sidor med sånt . 
Artiklar som skannades in för leverans och plötsligt försvann . 
Wow . Stal nån allt det där ? 
Du riskerar åtal för smuggling , skattebrott , och du hjälper inte dig själv . Du skrattar bort det som ett skämt . 
Jag vet inte vem som tog allt det där . Tänk efter . Jag säljer underkläder och munvatten och fotpuder . 
Saker som gör livet lite lättare för folk här uppe . 
Och vem vill ha kommunikationsutrustning ? 
Det har ingen praktisk användning . 
Såvida man inte vill sabotera Ranger . 
Dev Ayesa bröt strejken . 
Många är fortfarande förbannade för det . 
Kanske så förbannade att de bad dig om hjälp att hämnas . 
Varför skulle jag riskera allt ? Allt jag har byggt upp . 
Jag var mot strejken ända från början . 
Ni kan fråga vilka ni vill , de vet . 
Du vill att vi ber en hög terrorister att gå i god för dig . 
Nick Jennings var en god vän till mig . 
Visste du att hans dräkt smälte in i köttet ? 
Kan du föreställa dig vilken outhärdlig smärta han måste ha känt under sina sista ögonblick ? 
Jag hade inget med det att göra . 
Men för i ... - Hallå ! - Sätt dig , för fan . 
Hör på ! Ni bryter armarna av mig , för fan . 
Okej , så , du ska alltså ta dig genom åtkomsttunneln . Har du familj nere på jorden ? 
Ja . En bror och två systrar . Föräldrar . 
Det var ett tag sen vi ... Inte direkt ... Vad i helvete ? 
Kalla in alla . 
Vad fan ? 
Vad i helvete ? 
Vad i helvete ? 
