Albrightstipendiets kandidatträning 
Snabbare ! 
Hallå , San ! 
Ta det lugnt ! 
Skynda , Kwangmin ! 
Sakta ner ! 
- Herrn ! 
- Soldat . 
Varsågod . Bra jobbat . 
Herrn ! 
Varsågod . Bra jobbat . 
Tack , herrn . 
- Herrn ! 
- Soldat . 
Förlåt . 
Vad gör du ? 
Tar mat till min systerdotter , Jina . 
Du har mycket att tänka på . 
Det är okej . 
Oroa dig inte . Fokusera på studierna . 
Vad är bäst med utomlandsstudier ? Man slutar oroa sig för familjen och fokuserar på studierna . 
Jag ska göra det . 
Har din fars hälsa förbättrats ? 
Nej , han mår inte så bra . 
Jag ska bidra till dina levnadskostnader . 
Det behövs inte . Det är okej . 
Ta det . Jag insisterar . 
Tack , herrn . 
Då så , - ta din mat . - Okej . 
Uncle Samsik 
Uncle Samsik 
Far mot farbror 
Kang Seongmin gråter nog vid herr Ans fötter nu . 
Han vet inte att han svalde betet . 
Han är nog tacksam . 
Självklart är han det . 
Han har aldrig drömt om att bli premiärminister . 
Jag har haft honom runt lillfingret sen han var bebis . Vad gör alla amerikanska soldater ? 
Amerikanska soldater ? 
Nåt är på gång . 
De unga officerarna verkar hålla med om uttalandet . 
Amerikanska arméns högkvarter har ny information . 
Jag håller militären under kontroll . 
Vi kan muta nationalförsamlingen , men inte militären . 
Det såg vi under Japans ockupation . 
Vad för ny information ? 
Militären kan försöka ge förste infaterichefen makten . 
Förste infanterichefen ? 
General Choi Hanrim . Militären litar på honom och han står nära USA:s befälhavare . 
Choi Hanrim ? 
Kapitalförsvarsenhetens hemliga bunker 
Du träffade väl general Choi på Albrights avskedsceremoni ? 
Ja , det gjorde jag . 
Diskuterade ni statskuppen då ? 
Jag beundrade general Choi mer än nån annan i militären . 
Han hjälpte mig alltid . 
Han var som en far för mig . 
19 februari 1960 Seoul , Sydkorea 
Hotell Banya 
Honnör ! 
Kim San . 
Har du haft det bra ? 
Stämmer ryktet ? 
Jag gick med i demokraterna . 
Politik är ingen barnlek . 
Alla tror att de är annorlunda , men inser sen att de inte är det . 
Men då är det för sent . 
Jag ska minnas det , herrn . 
Ska vi ? 
General Choi respekteras av för många . 
Ska folk som respekteras bli beundrade ? 
Jag hatar dem . 
Där är han . 
Kim San står bredvid honom . 
Som sig bör . Det är hans mål i dag . 
General Choi är här . 
Står de inte varandra för nära ? 
Det är ju hans mål i dag . 
Det verkar ändå lite onödigt . 
Han är nästan Kim Sans fosterfar . 
En far heter Choo och en annan heter Choi . 
Hur många fäder har han ? 
Du är avundsjuk . 
Avundsjuk ? 
Å Cheongwooförbundets vägnar har An Kichul från Segangs Textilier nu donerat . 
I år skickar vi tolv stipendiater till USA . 
En applåd för Rachael Jeong från Albright . Min lillasyster . 
Damer och herrar . Rachael Jeong från Albright . 
Först och främst vill jag tacka er för er tid och jag uppskattar verkligen var och en av er här i dag . 
Vårt arbete är en ära . Men utan vidare dröjsmål är det mitt nöje att presentera Albrightstudenterna . 
Välkomna våra tolv stipendiater . 
Vi presenterar våra Albrightalumner . Kim San , Jeong Hanmin och Kim Kwangmin , kom fram . 
Givakt . Honnör . 
Rachael , har du pratat med ministern än ? 
Det var länge sen , överste . 
Vet din farbror ? 
När jag åker ... 
" Låt oss inte tröttna på att göra gott . Ty när tiden är inne får vi skörda om vi inte ger upp . " 
Galaterbrevet 6 : 9 . Ord jag lever efter . 
Så länge ingen av oss ger upp , kommer de frön vi har sått inte att gå till spillo . 
Du har inte berättat om mig ? 
Jag har inte berättat för min farbror , för han skulle bli besviken på dig . 
Överste , Albright har ögonen på dig och ditt tålamod . 
Om du börjar tröttna , ha lite tilltro . 
Tänk på vår kommande skörd . 
Jag ska hälsa min far och farbror . 
Ursäkta mig . 
- Farbror Samsik . 
- Michael . 
Min syster Rachael . 
Rachael , farbror Samsik . 
- Farbror Samsik . 
- Du vet väl vem han är ? 
Angenämt . 
Jag har hört så mycket om dig . 
Detsamma . 
Du låter som en amerikan . 
Jag är amerikan . 
Jag måste fixa mina skor . - Okej . 
- Ursäkta mig . 
Min sko ger mig problem . 
Vi ses . 
- Hej . 
- Hej . 
Cha Taemin stack efter att ha dödat tre av mina män . 
Slängde du alla bevis mot mig ? Det gjorde jag . Jag brände allt . 
Förresten ... 
Fortsätt . 
Under den senaste översvämningen sveptes en bro bort i min valkrets . 
Vi pratar om det sen . 
Visst . 
Jag sa det för att du gav mig klartecken . 
Ursäkta mig . 
Ja , fröken ? 
Kan du fixa min sko ? Jag ? 
Ska jag fixa din sko ? 
Ja , tack . 
Eller , glöm det . 
Jag löser det . 
Det är upp till dig . 
Ursäkta mig . 
Har du eld ? 
Minns du slaget vid Nakdongfloden ? 
Självklart minns jag . 
Vi bombarderades 28 timmar i sträck . 
Vad ska jag säga ? 
Jag trodde att du dog då . 
Ursäkta . Och jag tänkte för mig själv : 
" Vad gör kommunisterna här ? " 
Jag menar ... 
Vad är det ? 
Jag kan tolka åt dig om det går bra . 
Visst , det vore toppen . 
Jag undrade varför de inte skrattar åt mitt skämt . 
Ursäkta mig . 
Jag är hans tolk . 
Han ville säga : 
" Jag dog och kom tillbaka för att jag såg kommunister i himlen . " 
Det var ett skämt ! 
Jag berättade det . 
Jag trodde att jag var död . 
- Ja . - Ja . 
Han är rolig . 
Tänk att Kuba fick en kommunistisk regim . 
" Tänk att Kuba blev kommunistiskt . " 
Folk som du borde syssla med politik , general Choi . 
" Folk som du borde ... " 
Säg att det räcker . 
Det rör inrikesfrågor . 
Varför prata politik med en soldat ? 
Om Korea mot förmodan blir en kommunistisk stat ... 
" Prata inte politik med en soldat . " " Och om , jag säger om Sydkorea skulle bli ... " 
Jag tar över nu . 
Vem är du ? 
Jason Arrent ? Politisk tjänsteman på USA:s ambassad . 
Ambassaden ? 
Okej . Ambassaden . 
Varför lämnade du bordet ? 
Nån från ambassaden erbjöd sig att tolka . 
Du borde ha stannat där ändå . 
Vad pratade de om ? 
Ska han bli politiker ? 
Vad sa han ? 
Han sa : " Om Korea mot förmodan blir en kommunistisk stat ... " 
Ja , och ? 
Sen avbröt killen från ambassaden . 
Varför i ett så viktigt ögonblick ? 
Minns du mig ? 
Ja . 
Från stipendieceremonin . 
- Eller hur ? 
- Ja . 
Underbart . 
Du har bra minne . 
Jag minns allt från den dagen . 
Nationella rekonstruktionsprojektet . Det var intressant . 
En ögonöppnare . 
Tack . 
Tror du att det är möjligt ? 
Kanske . 
Om vi öppnar det , tar isär det och fixar det från grunden . 
Vad skrattar du åt ? 
Du fixade inte min sko . 
Du lät mig inte . 
Om jag gjorde det , hade du fixat den ? 
Många har förlorat pengar på investeringar i Kuba . 
Varför skulle nån vilja investera i Korea om det är ännu värre här ? 
Sydkorea är annorlunda än Kuba . 
Jag litar inte på Koreas regering än . 
Så ... Menar du att du inte tänker investera i vårt industrikomplex ? 
Vad mer behöver du ? 
Betalningsgaranti från Koreas regering . 
Betalningsgaranti ... 
Menar du allvar med att ge dig in i politiken ? 
Ja , herrn . 
Kan du stå upp mot vana politiker ? 
Jag ska göra mitt bästa . 
Kom och hälsa på snart . 
Jag vill diskutera nåt . Det ska jag . 
Du bugar mot hans bil . 
Vad sa Petron Harvest ? 
De bad om en betalningsgaranti . 
Det kan vi inte lova . 
Hoppa in . Låt mig skjutsa dig . 
- Hör av dig . 
- Vi ses . 
Bra jobbat . 
Lovade din kära fader Choi dig lite pengar vid sidan om ? 
Du är barnslig . 
Hur många fäder har du ? 
Färre än dina syskonbarn . 
Herregud . 
Så du har räknat dem ? 
Du borde lämna general Choi ifred . 
För att han är som en far ? 
Ska du döda honom också ? 
Vem tar du mig för ? 
Du erkände det själv . 
Du har rätt , det gjorde jag . Men ändå ... Det fanns omständigheter . Det var en sista utväg ... 
Att du lät Cha Taemin döda alla ? 
Jag ska få honom att lämna militären . 
Är det möjligt ? 
Jag har gjort det här hela livet . 
Vad är din plan ? 
Jag tar Pak Jiwook med Han Soo som lockbete . 
Och sen ? 
Sen tar jag Choi Hanrim med Pak Jiwook . 
Senaste nytt ! 
Kang Seongmin ambition bakom lokalt självstyre 
Senaste nytt ! 
Det kommer en artikel om ändringen av lokalt självstyre . 
Choi Minkyu kommer att tjata på Kang Seongmin om att få igenom den . 
Motståndare till ändringen tipsade media . 
Varför har du inte kontroll över partiet ? 
Få igenom den omedelbart . 
Men det tar tid ... 
Vi har knappt tid ! 
Gör vad som krävs . Sätt igång ! 
Vad sa han ? 
Han bad mig få igenom den . 
Direkt ? 
Är det möjligt ? 
Nationalförsamlingen 
Regeringen kan inte lägga sig i valet så öppet . 
Varför mobilisera regeringsarbetare inför valet ? 
Det är nödvändigt . 
Vi kan inte stödja en så orimlig ändring . 
Vi gör det för presidenten . 
Är du säker ? 
Inte för Kang Seongmin ? 
Mer än 20 års tjänst hos polisen lärde mig detta . 
" Alla har skelett i garderoben . " 
Ju närmare man tittar , desto fler skelett hittar man . 
Ni har förvaltat tillgångar under lånade namn , stört lokala företags anställningar , och mutat skolor att ta emot era barn . 
Jag har hämtat alla bevis från Nationella säkerhetsbyrån . 
Det som är bra för Kang Seongmin är bra för vårt parti , och i slutändan för presidenten . Okej ? 
Är Kang Seongmin med i Sineuialliansen ? 
Är det vad ni tror ? 
Kom ihåg att ni kan falla före honom ! 
Seonyoowon 
Jag samlade alla ledamöter som flydde till landsbygden . 
Det är bra . Vi kan få över 180 röster i morgon kväll . 
Lista på ledamöter som är för ändring av lokalt självstyre 
Förresten , det har skrivits fler artiklar . 
Jag tror att Samsik ligger bakom dem . 
Vem skulle Cha Taemin annars ha gett bevisen till ? 
Tipsade han tidningen om Sineuialliansen ? 
Låt oss prata om lagen om lokalt självstyre . 
Det är nåt skumt med Samsik . 
Jag skuggade honom . Han har umgåtts med Kim San , Choo Intaes svärson . 
De träffade An Yosub . 
Man kan inte lita på Samsik . 
Vem är Kim San ? 
Han jobbade på Nationella rekonstruktionsbyrån . 
Jag vill prata med dig , herrn . 
Han ser bekant ut . 
Har du inte läst tidningen ? 
Jag har träffat honom . 
Och ? 
Ska jag kolla upp honom ? 
Hallå ? 
Ja , han är här . 
Det är till dig , herrn . 
- Kang Seongmin . - Hej . 
Så det var där du var . 
Jag har nåt brådskande att diskutera . 
Vad säger du ? 
Ska jag komma över ? 
Visst , jag väntar . 
Vem var det ? 
Ta hand om ledamöterna från landsbygden . 
Vem var det , sa jag ? 
Var det Samsik ? 
- Den jäveln . 
- Jag tar hand om det . 
Du borde inte ... 
Du vet inte ens vad han kokar ihop . 
Jag tar hand om det . 
Var snäll och gå . 
Kära nån . 
- Starta bilen nu ! 
- Ja , herrn . 
Ta en titt . 
Meritförteckning Kim San 
Så herr An ersätter mig med Kim San ? 
Vilket är absurt . 
Det är otroligt . 
Misstänker han mig fortfarande ? 
Ska jag hålla ett öga på Kim San ? 
Om han visar sig vara ett hot , kan jag muta honom när det är dags . 
Tack . 
Ingen orsak . 
Jag gör bara mitt jobb . 
Även om alla sa åt mig att inte lita på dig , skulle jag ändå lita på dig . 
Vi måste driva igenom lagen om lokalt självstyre , va ? 
Ja , senast kl. 23.00 i morgon . 
Jag håller oppositionen på avstånd . 
Var försiktig . 
Du räddade mig när jag var i knipa . 
Jag ska göra även Yoon Palbongs del . 
Dags att gå hem . 
Vänta . 
Jag måste lätta på trycket . 
Nej , jag följer dig hem . 
Det är okej . Åk du . 
Bra jobbat . 
Säg åt Han Soo att samla alla . 
Taemin ? 
Sineuialliansen står upp mot den makt som förtrycker vårt folk . 
Sineuialliansen tyranniserar ingen för egen vinnings skull . " 
Taemin . " Vi motsätter oss allt och alla som monopoliserar makt och är beredda att använda våld och vapen . 
Alla som förespråkar förtryck ska straffas i Sineuialliansens namn . " 
Det är uppförandekoden du skapade när du var 16 år . 
Minns du den ? 
Den är Choi Minkyus verk . 
Jag skickade inte männen . 
Kang ... Seongmin är Sineuialliansens sista mål . 
Vänta . Ge mig en chans . 
- Att göra vad ? - Vad som helst . 
Jag gör allt . 
Vad som helst för att skärpa mig . 
Jag kan inte ... Jag kan inte dö så här . 
En chans ? 
Taemin , snälla ! 
En sista chans . 
Jag övervakar dig . 
Vad gör du här ? 
Vi måste prata . 
Följ med mig . 
Håller du kontakten med Yeojin ? 
Varför frågar du det ? 
Kang Seongmin agerar ut nu när han är trängd . 
Han vill ändra lokalt självstyre - och mobilisera ... - Är det därför du är här ? 
Det är offentligt . 
Varför är du efter honom ? 
Det sker en politisk reform efter valet . 
Ett parlamentariskt system införs och han blir premiärminister . 
Så du försöker stoppa honom ? 
Du ska få ett större scoop . 
Ett scoop ? 
En bild värd förstasidan på bråk i Nationalförsamlingen . 
Kang Seongmin vill få igenom lagen om lokalt självstyre . 
Det är din chans att etablera din närvaro . 
Ska jag ska gå emot honom ? 
Du lär dig snabbt . 
Vi vill få igenom lagförslaget så att han kan avancera i Liberala partiet . 
Jag har inget mer att lära dig . 
Genom att motsätta mig framstår jag som en kämpe för demokratin . 
24 februari 1960 Seoul , Sydkorea 
Nationalförsamlingen 
Är de liberala ledamöterna på väg ? 
Ja , även medlemmar utanför huvudstaden är på väg . 
Okej . 
Okej . 
Jag har samlat våra tio starkaste medlemmar . 
En har varit brottare . 
Vänta tills jag ringer dig . 
Okej . Men räcker tio ? 
Vi kommer att möta 100 personer . 
Du behöver inte oroa dig . 
Det går bra . 
Blockera dörren med dem . 
Vi går in . 
Lite dryck , tack . 
Här . 
Drycken är här . 
Varsågoda . 
Tack för er tid . 
Jag är nyfiken på Nationella rekonstruktionsprojektet . 
Tack för att du ska förklara det för oss oberoende ledamöter . 
Jag är Kim San , ekonomiutskottets ordförande . 
Angenämt . 
Ett nöje . 
Slå er ner . 
Vänta . 
Jag glömde viktiga dokument . 
Då börjar jag mötet . 
Bra . Jag kommer strax . 
Sätt er , allihop . 
Ledamot Sun , vad gör du här ? 
Jag glömde en sak . 
Hej , herrn . 
Ni är alla här . 
Kul att se er . 
Vi dricker lite te innan vi åker till Nationalförsamlingen . 
Det är inget speciellt . 
Jag vill bara tillbringa tid med er . 
Okej . 
Med tekniköverföringen från partnerbolag kan vår export överstiga en miljon dollar inom fem år . 
Borde inte ledamot Sun vara tillbaka ? 
Du har rätt . 
Han kommer säkert strax . 
- Vi går dit nu . - Ja . 
- Vad i ... 
- Vad har hänt ? 
Öppna porten ! 
Öppna porten , era jävlar ! 
Är ledamot Lee Chungwon här ? 
- Jag är här . 
- Där är du . 
Okej . 
Ska vi gå dit ? 
Inte än . 
Kom igen . 
Vi har varit här länge . 
Tänk att vi måste vänta så länge . 
Ge oss lite whisky . 
Ingen alkohol , sa han . 
Vem ? 
Samsik . 
Jag tar hand om det . Servera . 
Kom igen , var inte sån . 
Är ledamot Moon Kyungju här ? 
- Jag är här . - Okej . 
Ledamot Moon är här . 
Det är farligt , herrn . Snälla , kom ner . 
- Vem fan är du ? 
- Kom ner . Öppna dörren ! 
Hallå ! Öppna dörren nu ! 
Herregud . 
Mina herrar . 
Ni borde åka hem . 
Liberalerna röstar om ett lagförslag . 
- Nu ? 
- Vilket lagförslag ? 
Ändring av lokalt självstyre . 
Vi måste stoppa dem ! 
Vi fyra mot 100 ? 
Vad är vi , amiral Yi Sunsin ? 
Lagen om lokalt självstyre ? 
De försöker rigga valet ! 
Ledamot Kim ! 
Vad ska vi göra ? 
Vi har ingen chans . 
Vi borde ringa demokraterna . 
Jag ringer dem . 
Dags att åka till Nationalförsamlingen ! 
Åk till Nationalförsamlingen ! 
Skynda på ! 
Varför ska vi dit ? 
Kom igen . 
Kom igen . Skynda . 
Varför är ni kvar här ? 
Du kan inte stå rakt . 
Är det rätt läge för whisky ? 
- Jag går . 
- Senila dåre ! Tänk om Kim San blir skadad ? 
Gå ! Nu ! 
Vad är det med dig ? 
Hur vågar du ? 
Vad bad jag om ? 
Ska vi bara titta på ? 
Det är över 100 liberala ledamöter . 
Dags att rösta om ändringen av lokalt självstyre . 
Ni är väl inte här för att rösta emot ? 
Kom igen . 
Vi måste hindra dem . 
Vad sysslar ni med ? 
Hur vågar ni ? 
Vi knuffar oss in . 
Håll armkrok ! 
- Lagförslaget är ogiltigt ! 
- Det är ogiltigt ! Nej till illegala val ! 
Inga illegala val ! Lagförslaget är ogiltigt ! 
Vad i ... Släpp . Inga illegala val , Kang Seongmin . 
Hur vågar du attackera en ledamot ? 
Du är ingen ledamot . Du är Choi Minkyus lakej . Din lilla ... 
Herrn . 
Lagförslaget är ogiltigt ! 
Vi säger nej till illegala val ! 
Lagförslaget är ogiltigt ! 
Nej till regeringens inblandning i valet ! 
Säg nej till illegala val ! 
Lagförslaget är ogiltigt ! 
Vem gjorde så mot ditt stiliga ansikte ? 
Vem annars ? 
Kang Seongmin . 
Bra jobbat . 
Jag gör det . 
Oroar Kang Seongmin dig ? 
Självklart inte . 
Du verkar ha varit med och drivit igenom lagändringen . 
Ska vi prata om valfusket ? 
Får jag röka först ? 
