TIDIGARE ... 
Morfar ? 
- Vad gör ni ? 
- Inget . 
Det går ändå inte att se Saturnus . 
Tänk om någon ser vagnen gunga och tittar in ? 
Vi hittade Van , han är på ett flyktingläger i Malaysia . 
Jag känner en malaysisk man . 
Han kan tänkas hjälpa er , men han tar betalt . 
Helsike . 
Jag behöver en läkare . 
- Känner du någon ? 
- Det är klart . 
Jag tror att jag är gravid . 
De brydde sig inte om oss när de utsatte oss för radioaktivt nedfall med de där testen . 
Jag har aldrig pratat om det , och tänker inte börja nu . 
Jag vet inte vad jag ska göra med Mia . 
- Vad skulle du göra annorlunda ? 
- Inget . 
Du är perfekt . 
Jag vet att du kan fixa den . 
Största hedersmärket som jag har sett . 
Min bräda , jag åker först . 
Morfar . 
Snälla , hjälp ! 
Snälla ! 
Ingen pacemaker ? 
Klockan . Jag vet inte om den är uppdragbar eller batteridriven . 
Den har stannat . 
Uppdragbar . 
Då sätter vi den tillbaka . 
- Är du säker ? 
- Det är klart . 
Nej . 
Du kan lämna ringen . 
Mormor ? 
Vita . 
De begraver sina döda för snabbt . 
- Hjälp mig att förstå . 
- Kröningskyckling . 
Det är morfars favorit sedan drottningen kröntes . 
Jag tycker vi borde skicka dem tillbaka till drottningen . 
Vet du vad ? Jag har funderat . 
Kanske vi borde skicka pappas aska tillbaka till England . 
- Ölen är inte kall . 
- Ja , det är så han gillade den . 
Mamma frågade just vad vi borde göra med morfar . 
Skicka honom till London , kanske ? 
Skjuta ut honom ur en kanon ? Jag vet inte . 
Skaffa en gravplats här ? 
Ja , kanske vi borde ha en här och en i Storbritannien . 
Eller något däremellan ? 
- Som till havs ? 
- Okej . 
Mia kunde göra det på sin bräda . 
Det är en bra idé . 
Pappa älskade havet . 
Nej , ingen chans . Inte jag . 
Jude . 
Hur klarar du dig ? 
Jag är okej . 
Han ... 
Bob , han ... 
Han levde ett gott liv . 
Men efter att mamma dog , hade han aldrig någon annan . 
Det hade varit trevligt om han hade hittat kärleken igen . 
Ursäkta mig , Eileen . 
Kan du ta hand om de här ? 
Jag för ut de här . 
Jag tog med en vän . 
Minns du " Sam " ? 
Sambuca . 
Det tar tid att smälta . Sorg . 
När jag miste Frank , trodde jag smärtan aldrig skulle ta slut . 
- Det blir bättre , eller hur ? 
- Inte egentligen . 
Vi slapp tänka på jobbet åtminstone . 
Inte jag . Jag är fortfarande besatt . 
Vad fan är det Wayne planerar ? 
Envis som han är , dum som han är , vem vet . 
Är det här som festen är ? 
Låt mig presentera dig för min svåger , Mick . 
Han är familjens entreprenör . 
Trevligt att träffas , mr Entreprenör . 
Jag försökte få det att funka med Tony . 
- Men du vet säkert hur det var . 
- Jag avskedade ju honom först . 
Ska du gå nu ? 
- Ja , min skjuts väntar . 
- Russell ? 
Varför bjöd du inte in honom ? 
Du vet att han är välkommen . 
Av dig . 
Du vet om din grej , va ? 
När alla känner sig vilse , gör du din grej . Du tar kontroll . 
- Gå din väg . 
- Så är det . 
Missförstå mig inte , din familj är toppen , men fan vad jag hatar folkmassor och uniformer . 
Du passar i kostym . 
Åh , sluta . Jag kvävs . 
- Okej , vi ses . 
- Nej . Inte än . 
- Jag är inte färdig med dig . 
- Jag måste gå . 
Här har du den . 
Vinner inga skönhetstävlingar . 
Tack , Spindeln . 
Efter det här ska vi surfa . 
Inte nu . Inte än . 
Du ska inte vänta för länge . 
Först är det en vecka , sedan månader . 
Plötsligt har det gått ett år . 
Nästa gång du ser en stor våg där ute , ska du ta dig dit . Okej ? Bara andas , och surfa . 
Fint av Bob att fixa din bräda , men det behövde inte göras . 
Som jag sa , det är ett hedersmärke . 
Gå . 
- Gamle Bob , va ? 
- Gazza . 
En påminnelse om att ingen undgår liemannen . 
Min svärfar måste alltså kola av innan du skulle dyka upp . 
Hej , det är stängt . Privattillställning . 
Jag vet . 
Jag är här två dagar till , om vi inte pratar ... 
- Det här gjorde de mot oss . 
- Han ska just gå . 
Dags att gå , kompis . 
Har du inte berättat för henne ? 
Lyssna , George . 
Helvete . 
Om du inte är sjuk än , är du skyldig oss det . 
- Är du okej ? 
Låt bli , Tony . - Hallå . 
Varmt öl och engelska mackor var inte så populärt . 
Vad handlade den där scenen om ? 
Du anföll en sjuk man inför familj och vänner . 
Han sa saker om Bob . 
Jag knuffade honom inte , han föll . 
Som vad ? 
Jag vet inte . Men han sa att Bob var skyldig honom pengar . Han ville ha pengar . 
Han verkade känna dig , inte pappa . 
Han talade skit om Bob , och jag blev arg , okej ? 
Älskling , vad är det ? 
Jag sa ju . Ingenting . 
Okej . 
- Vart går du ? 
- Till kontoret . 
Miss Kulkova , ursäkta att ni fick vänta . 
Labbet är långsamt den här tiden på kvällen . 
Du är alltså gravid . 
Fantastiskt . 
Grattis . 
Ungefär 16 veckor . 
Du är i god form . 
Tack . 
Vi är väldigt glada . 
Bra . 
Jag måste låsa här , ni hittar säkert ut själva . 
Vi ses om sex veckor . 
- Tack så mycket . 
- För all del . 
Yvgeny , funktionärerna . 
Ingen vill det här . 
Vad vill du ? 
Vad jag vill ? 
Det kvittar . 
En gravid miss Sovjetunionen skulle skämma ut hela landet . 
Och pappan ? 
Han är en skit . 
Har du sett mina kläder ? De där klänningarna . De syddes till mig för länge sedan . 
Jag ryms inte i dem , de skickar hem mig . 
Vi hittar på något . 
Jag behöver en drink . 
Du också ? 
Sådant oväsen . 
Vi går och lägger oss . 
Jag behöver bara en stund . 
Kom igen , Bob . 
Låt mig sova lite . 
Han hatade de här kungliga smörgåsarna . 
Du ser trött ut , mormor . 
Ja . Tack vare Bob . 
Han gillar dig fortfarande . 
Du vet vad du måste göra . 
Doris kan hjälpa . 
Ja . Jag vet . 
Din middag är klar om två minuter . 
Säg till din pappa att du fick extra musslor . 
Tack , mr Mui . 
Du har fullt upp . 
Vi är gasdrivna . 
Ingen strejk stoppar oss ! 
Hemuppgifter ? 
Jono sa att du var professor . 
- Ingenjörsvetenskap . - Jaså ? 
Jag försöker räkna ut var Skylab kommer att störta . 
Kan du ta en titt på det ? 
Varför ett fysikproblem ? 
Det är ett fysikproblem . 
Varför inte en linjär regression ? 
Troi oi . 
Lyssna inte på honom . 
Han tror allt är en linjär regression ! 
Lam , var är kaffeskeden ? " Linjär regression ! " 
Han ställer alltid till problem . 
Carl Friedrich Gauss tittade på himlen . 
Han visste det fanns en annan planet , fast ingen hade sett den . 
Han hade ingen räknare . 
Det är inte matematik . Det är statistik . 
Hur gör jag det med Skylab ? 
Nu ... 
X , Y. Börja enkelt . Bara två dimensioner . 
Är det öppet ? 
Ja , alltid öppet . 
Ingen går hungrig , min vän . 
- Hej . 
Svetlana ? 
- Hon är upptagen . 
Jag har just gått sex trappor upp . 
Vi är bekymrade över Svetlanas figur . 
Hennes vikt . 
Det är garderobsavdelningens problem . 
Vad ville hon ? 
Det västerländska livet gör dig mjuk . 
Om du förlorar , är det illa för oss . 
- Vad ? 
- Du äter vad jag säger . 
Motionerar när jag säger . 
Nej , nej . Vi måste bara hålla Lydia nöjd . 
Jag tar hand om henne . 
Men vi måste sköta det bra . 
De tittar på oss där hemma , eller hur ? 
Hjälp mig vinna henne på min sida . 
Det är inte en skönhetstävling . Det är en popularitetstävling . 
På akademin var jag bäst på tvångsåtgärder vid förhör . 
Nej . Skräm henne inte . Bara charma henne . 
Jag bjuder henne på lunch . 
Jag flörtar med henne , hon gillar det . 
Du vinner och får en hjältemedalj . 
Jag åker hem och Niki kommer tillbaka . 
Nu måste jag hitta Bobs " malaysiske man " . 
Han känner någon på flyktinglägret . 
Bob gav honom våra pengar . Han är i Bayswater . 
Bayswater ! Mr Teo ? 
Mr Teo ? 
Han har ett brett leende , han ser omtänksam ut . Som de som råder att föda upp vaktlar . Han lovar dig världen . 
Vet du var han är ? 
Han är lögnare . En skurk . Säger vad som helst för att få dina pengar . 
Han säger alltid , " Jag jobbar på det , lah . " Ber du om dina pengar , hotar han anmäla dig . 
Ursäkta . 
Är du okej , em ? 
För att minimera fel , tar man förstaderivatan och sätter den till noll ? 
Minimera inte fel ! 
Positiva och negativa stryker ut varandra . 
Kvadrera residualen . Ser du ? 
Saknar du inte att vara professor ? 
Jag miste mycket mer än bara mitt jobb . 
Ja , min kaffesked ! 
Här har du din sked . 
Men för att räkna behöver du data . 
Trettio observationer , annars går det inte . 
- Tror du att det räcker ? 
Okej . 
- Börja där . 
- Trettio ... 
Du är inte den tuffing som du ser ut att vara . 
Du bryr dig om dessa flickor som om de vore dina döttrar . 
Min första kommendant . 
Han lät oss stå ute på vintern . 
I Sibirien . 
Inga handskar . 
Fick man en köldskada , avlägsnade han fingret själv . 
Personligen älskar du dessa flickor så . 
Har du döttrar ? En fru ? 
Min fru ? 
Cancer . 
Jag har en son , Nikita . 
Niki . 
- I armén . 
- Livet är hårt där , va ? 
Livet kan vara hårt var som helst . Visst ? 
Men vi vet hur man dricker . 
Som före detta miss Adelaide , vet jag hur man böjer på armbågen . 
" Böjer på armbågen ? " 
Särskilt med en snygg utländsk agent . 
Så Svetlana kommer att vinna , va ? 
Miss Universum har standarder . 
Svetlana måste ta hand om sin vikt . 
Annars låter jag inte henne gå på scenen . 
Jag tar hand om Svetlana . 
Det är inga problem . 
Låt oss " böja på armbågen " . 
Hej , du har ringt Lawley familjeplaneringsmottagning . Vi kan tyvärr inte ta ditt samtal ... 
Kamrat . Vi har ett problem . 
Det är dags , Nan . 
Inte än . 
Är du redo , Eileen ? 
Okej . 
Vi ses , Bob . 
Vi ses på andra sidan . 
Trevlig doft ? 
Vi hjälper din pappa gå vidare . 
Han har besökt mormor i flera dagar . 
Besökt Eileen ? 
Ja . 
- Skylab kommer att krascha här ! 
- Är det på nyheterna ? 
- Linjär regression . 
Lam visade mig . 
- Har han fortfarande öppet ? 
Ja . Han behöver inte er . 
- Han har mer jobb än någonsin . 
- Lams mat är jättegod men du måste rådfråga experter . 
- Hur är det med CSIRO , NASA ... 
- Vi gjorde beräkningarna , mamma ! 
Bara en liten bit kan förstöra vårt hus . 
Ibland händer det hemska saker , Tilly . 
Och ... Beräkningar kan inte ändra på det . 
- Pappa ! Skylab kommer att krascha här ! - Vad ? 
Tilly ... 
Vi måste berätta för alla . 
CSIRO . Alla ! 
Hon är precis som du . 
Som sprider nyheter om undergång och olycka ? 
- Jude ... 
- Jag menar , jag har ... Vi har varit utan el i flera dagar . 
Jag har försökt allt . 
Jag tar fortfarande hand om pappas saker . Och sen ... 
Låt mig fixa det här . 
Varför tar du inte paus ? 
För att jag är okej . 
Jag är okej . 
Judy . 
Du är den enda som inte har tagit tid att sörja . 
Vem var mannen på vakan ? 
Jude , jag var en idiot , okej ? 
Jag är ledsen . 
Förlåt . 
Tony , varför berättar du inte för mig ? 
Vad är det som pågår ? På riktigt . 
Det som pågår är att jag letar efter stearinljus , så att ficklampan inte dör , okej ? 
Jude ... 
STREJKBRYTANDE BITCH BRYTER 
Det är tidigt . 
- Ja . Bärgningsbilen kommer idag . 
- Nej , du kan inte göra dig av med den här . 
- Mia ... 
- Nej . Allt kan inte gå idag . 
Husvagnen , hans aska . 
Mia . 
Jag är ledsen , mamma . 
Jag vet att morfar skulle ha velat det , men jag tror inte att jag kan . 
Älskling , ingen ber dig göra det . 
Jag tror inte att jag är redo . 
Vet du vad ? 
Jag tror den här tillhör dig . 
Jag frågade morfar en gång , om han någonsin tänkte hur det hade varit , om vi inte hade åkt från England . 
Vet du vad han sa ? 
" Aldrig . 
Jag skulle frysa tuttarna av mig . " 
Det sa han . 
Och ... " Vi skulle inte ha någon Mia . " 
Kanske jag borde . 
Men husvagnen stannar . 
Mitt arv . 
Och hans gamla handduk , den behåller jag . 
Eileen . 
Eileen . 
Vi har en grej för pappa på eftermiddagen . 
Bara för de allra närmaste . 
Okej . 
Jag vore glad om du kom . 
Du borde vara där . 
- Jag vill inte ... - Jude . 
Tack . 
Tack för att du älskade honom . 
Vi kunde ha firat jularna ihop . 
Jag ville berätta för dig . 
Det skulle inte vara en hemlighet . 
Du behöver inte förklara . 
Jag visste inte vad vi var tills nu . 
Och nu är det för sent . 
PRODUCENTERNA TACKAR RESPEKTFULLT ABORIGINERNA OCH FOLKET PÅ TORRES STRAIT-ÖARNA DE SOM ENLIGT TRADITION ÄGER MARKEN OCH HAVET DÄR DETTA PROGRAM SPELATS IN 
SKAPARNA VILL BEAKTA NOONGARFOLKET . RÖKRITER ÄR VIKTIGA I KULTUREN . 
PYRANDE VÄXTERS RÖK RENAR EN PLATS OCH PERSONERS ANDE , KROPP OCH SJÄL . 
