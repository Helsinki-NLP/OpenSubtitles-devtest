Ordning i rättssalen ! 
Åklagare , fortsätt . 
Jag frågar en gång till . 
Under uppdraget såg du den tilltalade döda civila eller inte ? 
Svara på frågan ! 
Ska du inte svara ? Är det mamma ? 
Vem är det ? 
Det är Juncheol . 
Vem gav dig numret ? 
Det är inte viktigt . 
Bale lever fortfarande . 
Han är på väg till din mammas begravning med Seongjo Lee . 
Snälla , svara ! Kom igen ! 
Vad i helvete ? 
Ursäkta , min telefon dog . 
Får jag låna din och ringa försäkringsbolaget ? 
Helvete ! 
Släck lampan ! 
Vad fan ? 
Så spännande . 
Våning två i mitten ! 
Eldupphör ! 
Hur går det ? 
Helvete . 
Kom in . 
Hör du mig ? 
Hallå ... 
Vad fan ? 
Det är inte din turdag idag . 
Må du finna inre frid . 
Vad fan händer ? 
Är alla döda ? 
Allt var serverat på ett fat . 
För guds skull . 
Vad tar er så lång tid ? 
Kan ni skynda på ? 
Skjut mot taket ! 
Du skulle ha säkrat din sikt i mörkret . 
Du har förlorat din skicklighet . 
Minhye . Nån som du är värd att ta med till helvetet . 
Åh ... Hej , Jian Jeong . 
Jag är Bror . 
Sätt på de där . Sätt dem på Jeongmin . 
Va ? 
Hur vet du vem jag är ? 
Va ? 
Jag kan snurra den hela kvällen . 
Dessa sex har hyrt åkturen . 
Ni måste vara rika . 
Tjejen som blundar och killen i skinnjackan . Är ni släkt ? - Eller ett par ? - Håll i mig . Va ? Håller ni hand ? 
Titta på det där . 
Jag tillåter det inte . Attack ! 
Vad händer nu ? 
Sitt inte där . 
- Förklara dig ! - Junmyeon . Rör dig inte . 
Då ramlar du igen . 
Tjejen har de starkaste benen jag någonsin sett ! 
Titta så hon kniper ! 
Tack . 
Då går jag in då ... 
Jian . 
Kan du inte vänta ? 
Va ? 
Ska jag göra något innan jag går in ? 
Du har ingen koll alls , va ? 
Jag lagar den för 50 000 won . 
Här är min farbror . 
Jaha ... Hej . 
Du är för ung , kör utan hjälm och med olagliga modifieringar . 
Visa körkortet . 
Lägg av . 
Du är så gammalmodig . 
Låt ungdomarna pussas . 
Jian , så här . 
Jag vill se ändå . 
Visa ditt körkort . 
Jag har det inte på mig . 
Jag borde åka . 
Trevlig kväll . 
Jag följer med dig . 
- Jag ringer dig ! 
- Kom här . 
Va ? Ska du med ? 
Kör till affären . 
Såg du att han inte bugade när han hälsade på mig ? 
En bulgogiburgare och två räkburgare . 
Hon har jobbat här ett tag . 
Hon jobbar på gimbap-stället också . 
Bor hon hos sin farbror ? 
Farbror , älskare , hallick , vem vet ... 
Det är hennes farbror . 
- Ja . - Så känslig . - Så känslig . 
- Inte alls ! 
- Du är hemsk . - Hon är sån . 
Varför ? 
Inga föräldrar ? 
Just det , du vet inte ... Du började hos oss sent . 
Hör på . 
Hennes mamma och pappa ... Vill du bli slagen med 
- en stol igen ? - Traumat ! 
Smaklig måltid . 
Minsook , umgås ni ? 
Kom , vi går . - Va ? - Varför ? 
- Vi går . - Varför ? - Va ? - Nu går vi . Kom . 
- Vad ? - Bara ... 
- Vem är hon ? 
- Ingen . 
De har beslagtagit fyrahundra vapen , fem armborst och trettiotvå elpistoler . 
Den som ertappas med att bära vapen utan tillstånd riskerar upp till 15 års fängelse . 
Du var konstig mot Minsook . 
På mellanstadiet när hon var hemma hos oss ... 
Du stirrade på henne i tio minuter som ett pervo . 
Det kostade mig min enda vän . 
Och Jinki , privatläraren . 
Han skojade bara lite . Du hotade honom , och dagen efter slutade han . 
Hör på , Jian . 
För det första , Minsook stal min klocka den dagen . 
Jag tittade på henne för att bekräfta det . 
Hon lämnade tillbaka klockan efter . Och så var det med det . 
För det andra , privatläraren , Jinki ... 
Han greps för ofredande veckan efter . 
Det är mitt jobb att skydda dig . Jag gjorde mitt bästa . 
Junmyeon då ? 
Vad gjorde han ? 
Man får inte köra motorcykel så ung . 
Och utan hjälm ! 
Och han röker ! 
Han stank av rök . 
Lägg av ! 
Farbror . Vet du varför jag har två jobb ? 
För att ha råd att flytta härifrån . 
Jag har funderat på varför jag inte är som alla andra . 
Du uppfostrade mig , men ... Försöker du hålla mig inlåst ? 
Jag är ingen mönsterelev . Men jag är inget problembarn heller . 
Varför lägger du dig i allt ? 
Jag vill umgås med vänner som alla andra . 
Och jag vill dejta . 
Får jag det ? 
Om du kan göra en sak ... 
I ansiktet . Slå mig en gång , så får du flytta . 
Jag menar allvar . 
Jag med . 
Är du klar ? 
Jag dukar av . 
Döljer du något för mig ? 
Mamma och pappa ... Dog de på det sätt som de säger ? 
Jag minns faktiskt inte . 
Du måste berätta . 
Tänker du slå mig ? 
Det var svårt att ta upp det här ! 
Vad är det ? 
Du undviker frågan . 
Glöm det och bo kvar då . 
Du är så långsam . 
Du får diska . 
Du är så irriterande ! 
Sväng höger . 
Så där ja . 
Lite till . 
Bra jobbat , Jian . 
Långsamt . 
Hissa ner mig . 
Okej ! 
Wow , Jian ! 
Du klarade det . 
Du är duktig ! 
Bra jobbat . 
Parkera den , sen äter vi . 
Flytta på dig ! 
Flytta på dig , sa jag ! 
Flytta på dig ! 
Vad gör du , Jian ? 
Du skrämmer mig ! 
Bara subbor bråkar med sin familj . 
Lägg dig inte i , Pasin ! 
Fällde du mig ? 
Du är långsam som en snigel . 
Du kan inte röra honom . Inte ens nudda . 
Varför är ni på mig ? 
Släpp mig ! 
Släpp mig ! 
Släpp mig ! 
Hallå ! Släpp mig ! 
Släpp ... 
Du har gjort fel . 
Hur kan du göra fel varenda gång ? 
Du är så irriterande . 
Jag tog ut den ! 
Titta . Fel igen . Hur kan du mäta fel varenda gång ? 
Sluta gnälla . 
Svimmade jag ? 
Jian är vaken . 
Du måste ha varit jättetrött . 
Svimmade jag ? 
Hur kunde du låta din niece svimma ? 
- Va ? 
- Hon har rätt . 
Det var han ! Inte jag . Ja . Va ? 
Du sa åt mig att göra det . 
När då ? 
Vilken lögnare ! 
Fan ta dig ... Gå och dö ! 
Du sa åt mig att göra det . Du tvingade mig . 
Otroligt . När då ? 
Parkera gaffeltrucken ! 
Vad har du för hand ? 
Hit med huvudet . 
Förlorare får stryk . 
Lodisar . Betala först . 
Okej . 
Pasin , det du gjorde mot mig tidigare ... Lär mig . 
Ska jag lära dig thaiboxning så att du kan slå Jinman ? 
Ja . 
Nej . 
Ja , mästare . 
Smyg fram och slå honom när han sover . 
Men är inte det att fuska ? 
Det verkar för lätt . 
Tror du det ? 
Jag vill flytta hemifrån . 
Jag kan inte bo med honom . 
Den thaiboxning som jag tränar är tuff . 
Du klarar det inte . 
Jo . 
Jag gör allt du ber mig om . 
Tre gånger i veckan . 500 000 won i månaden . 
Jag har inte så mycket pengar . 
Jian . Jag måste skicka min son till privatskola nästa år . 
Så jag behöver mycket pengar , men jag har inga . 
Jag borde bara dö . 
Jag tjänar inte mer än 50 000 won i veckan . 
Taget . 
Följ mig . 
Lektion ett . 
Börjar vi nu ? 
Blockera mig . 
Ett , två . - Ett , två . - Armbågarna upp . 
Bibehåll formen . 
Håll balansen . 
Jian ? 
Du är för stel . 
Är du bättre ? 
Det var på öret . 
Ett , två . 
Snigel . 
Snigel , du är så långsam ! 
Res dig upp , Snigel . 
Hej ! 
Vad gör du ? 
- Sätt ner mig . - Så långsam , Snigel . 
- Skynda ... - Jian ? 
Vad i helvete ? 
Du är söt . 
Vilka var de ? Dina vänner ? 
Vi är bättre . 
Skrämde vi dig ? 
Du är väldigt vacker . 
- Visa ditt ansikte . - Minsook ? 
- Du . - Jian ! 
- Du ! - Vad fan ? Vad i helvete ? 
- Helvete . - Vem fan är du ? 
Du förstörde allt ! 
Salladslök ? Är det här ett jävla skämt ? 
Bra . Jag är sugen på ramyeon . 
Du ... Hon stack , så du får gottgöra det . 
Kan du det ? 
Jävlar . 
Vem fan pratar jag med ? 
Vad glor du på ? 
Vad är det ? Vad försöker du göra ? 
Är du en boxare eller något ? 
Vad är det ? Vill du leka ? 
Vad i ... 
Du är ny här . Det räcker . 
Hör på , Jian . 
Jag vet att Pasin har gjort dig starkare , men det räcker inte mot någon med kniv . 
Spring nästa gång . 
Släpp av mig hos Pasin . 
Jag behöver mina 350 000 won för att betala hyran ! 
Han är borta sen tre dagar . 
- Han stal 500 000 won . - Lugna ner er . 
Vi ska kolla allt . - Vänta bara . - Vad är det som pågår ? 
Jian ! Pasin , den jäveln ! 
Han lånade pengar och stack . 
- Va ? - Inte bara mina ! Alla här lånade honom pengar . 
Vad ska vi göra ? Vi är körda ! 
Är Jian Jeong här ? 
Det är jag . 
Jian , du är ingen snigel längre . 
Vad är det här ? 
Är det din skola ? 
Det finns en i badrummet . 
Du är galen ! 
Hur länge har du tittat på mig ? 
Vem byggde detta ? 
Min farbror ? 
Inte nu , Jian . 
Minhye har slut på kulor . 
Fler män kommer snart ! 
Det slutar inte här . Chefen sa det ! 
Minhye får inte dö om vi vill stoppa dem . 
Vi måste ut dit och ge henne fler kulor och medicin ! 
Vad i helvete säger du ? 
Vänta ... Det är för ljust ! 
Det är för ljust ! 
Xeroderma pigmentosum . Xeroderma pigmen ... 
Om jag ... Om jag utsätts för ljus länge gör det ont ! 
Släck ljuset ... 
Skynda ! Släck ljuset ! 
Du har inte svarat än ! 
Vad är allt detta ? 
Hur länge har du iakttagit mig ? 
Du kom till det här huset den 26 juni 2009 . 
Jag kom till det här huset den 20 juni 2009 . 
På bara ... 
Så där ja . 
Han spelar bara för att väcka sympati . 
Vad gör han här ? Han spionerade på dig . 
Jag ska sätta mig in i varuhusets system . Vi kan få veta mer om din farbror . 
Vad är det här ? 
Varför har ett vapenvaruhus ett sånt här serverrum ? 
Jian ! 
Lita inte på honom ! 
Öppna ! 
Vad gör jag nu ? 
Nej . 
Släpp mig . 
Släpp mig , skitstövel . 
Jian Jeong ? 
Öppna den andra lådan till höger . 
Ett . 
Om ägaren av murthehelp , Jeong Jinman , dör eller är frånvarande , ärver Jeong Jinmans niece , Jeong Jian , murthehelp . Två . När Jeong Jian tar över murthehelp kommer hon att samarbeta lojalt och sköta uppgifter som redovisning , ledning och personalhantering . 
Tre . Vid överlämnandet har Jian Jeong rätt att avstå från sitt arv ... 
Hon bekräftar med signatur ... Sex . Om överlämnandet sker enligt dessa regler ... Nödvändiga åtgärder vidtas ... 
Tio . Som murthehelp-anställd lovar jag att följa murthehelps ägares order , vad de än må vara . Och jag ska riskera mitt liv om så krävs . 
Jag läste allt . 
Berätta nu om du samtycker till att ta över murthehelp . 
Det finns papper och penna . 
Chefen planerade allt . 
Han räknade med att dö och att murthehelp skulle attackeras . 
Följ nu bara min guide ... 
Släpp Jeongmin , nu . 
Nej . 
Jag kan inte . 
Du skulle ju lyda mig . 
Du lovade . 
Minns du inte ? 
Släpp Jeongmin nu . 
Vad som helst , men inte det . 
Det finns ett skäl . 
Vad ? 
Jeongmin orsakade chefens död . 
Jeongmin ! 
Sluta . 
Vad gör du , Jian ? 
Tror du verkligen på honom ? 
Håll käften ! 
Nej . 
Nej , Jian . 
Jian . 
Tänk efter . 
Jag var med dig när vi nästan dog nyss . 
Och en kvinna drogade mig . 
Minns du inte ? 
Jag hjälpte till med webbplatsen och begravningen ! Skulle jag ha dödat honom ? 
Du undanröjde nog bevis under begravningen . 
Undanröjde vad ? 
Jag hittade hans telefon , och på grund av det hände allt , och jag dog nästan ! 
Jian . Han då ? 
Vet vi ens varför han är här ? 
Har han bott under er hela tiden ? 
Är det normalt ? 
Är han en parasit eller ? 
Jian Jeong . 
Är det inte konstigt att ... 
Håll käften ! 
Du tittade på Jian naken , pervo ! 
Nej ! 
Din farbror skulle aldrig begå självmord . 
Jian . 
- Lyssna inte ... - Tyst ! 
Jag vill höra hans version . 
Självklart . Visst , Jian . 
Men tänk efter noga . 
Det här är löjligt och orättvist . 
Fortsätt . 
Han kom till chefen . Sen dog chefen . 
Om du är nyfiken , öppna videon märkt " 0404 " på skärmen där borta . 
Du ... Vad gör du ? 
Är du en hacker ? 
Nej ! 
Nej , klicka inte på den . 
Vi vet inte vad som händer om du gör det . 
Dörrarna kan desarmeras så att mördarna kan komma in . 
Se dig omkring . 
Nej . 
Skynda dig , klicka på den . Titta på den . 
Han kanske ligger bakom allt . 
Nej ! Det är inte sant ! 
Han ljuger ! Klicka på den nu ! 
Jian ... Vänta , Jian ... 
Minns du ? Den som berättade för din farbror att du var inlåst i skolförrådet var jag . 
Här . 
Här ! 
Hör på , Jian . 
Beslutet är helt och hållet ditt . 
Vad ska du göra ? 
Behålla eller ge bort den ? 
Behålla den . 
Jag har döpt honom . 
Dooney . 
Jag ska ta hand om Dooney . 
Okej . Gör så . 
Men ... Hör på , Jian . 
Alla val du gör kommer med ansvar . 
Om Dooney dör , måste du ta ansvar för din sorg också . 
Du får gå . Ge kvinnan vapen och medicin . 
Okej . 
Det här är en present . 
Kan du ge mig mössan ? 
Just det ... 
Lämna inte varuhuset , vad som än händer . 
Lova ! 
Gör det inte . 
Vem är du ? 
Minhye . Det är jag . 
Det var längesedan . 
Du har växt . 
Mår du bra ? 
Jian . Tack . 
Tack för att du valde mig . 
Ja , visst ... 
Men ... Visste du ? 
När vi var små ... Den som låste förrådet var jag . 
Vad var det ? 
Samma som jag fick . 
Det fungerar bra . 
Dooney ... 
Du ... Vem är du ? 
Hur fungerar den ? 
Har den en knapp ? Inte mer ? En , två , tre . 
Jäklar ! 
Styr du den med datorn ? 
