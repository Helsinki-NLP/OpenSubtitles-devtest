TIDIGARE I SERIEN ... 
- Gazza kastade den . - Vad ? 
- Han skulle aldrig göra det . - Men det gjorde han . 
Har du varit här i några år ? Och Vietnam , bara lämnade du . 
Du hjälper mig att hoppa av . 
Skylab kommer att störta här . 
- Sades det på nyheterna ? 
- Linjär regression , Lam visade mig . 
Tack för det här , pappa . 
Vi gör vad vi måste göra , för att vara trygga . 
Håll det kort och sött . Med betoning på " sött " . 
Du är beviset på hur långt aboriginer har kommit under de senaste 150 åren . 
Säg mig , Eileen , hur många av dessa år har du bott i Scarborough ? 
Det sades till mig nyligen att jag aldrig ska glömma mitt förflutna . 
När jag var ung bodde jag på min makes marker , tills vi blev fösta till Yalata Mission för att bana väg för brittiska och australiska regeringens kärnvapentest . 
Du kanske känner till platsen . 
Maralinga . 
DOULL STRÖMFÖRSÖRJNING Är du okej ? Säkert ? 
Tänker du lära dig japanska medan du syr balklänningar ? 
Jag måste få veta vad Waynes papper handlar om . 
- Du är galen . 
- Märkte du det först nu ? 
Klänningarna kanske gör slut på mig . 
Men strejken gör det inte . 
Så ska det låta . 
Vi fixar skiten . 
Bara inget händer under Miss Universum-sändningen . 
Eller mot rymdforskarna som varnar oss för Skylab . 
Åtminstone behöver vi inte genomleva konsekvenserna . 
Apokalyps är ett sjujäkla sätt att sluta en strejk på . Men pluggisarna säger att Skylab landar i Indiska oceanen . 
En exploderande rymdfarkost ? 
Det hade varit för lätt . 
Gazza ? 
Någon jävel skar sönder mina däck . 
Behöver du skjuts ? 
Tack , men ... Jag är okej . 
Kom igen , Gazza , hoppa in . 
Jag kör hem dig . 
Hur mår du ? 
Bra . Jag mår bra . 
Jag lyssnade på den här när tegelstenen träffade vindrutan . 
Den som kastade den förstörde också sången för mig ! 
Mitt livs mest skrämmande ögonblick . 
Jag förstod inte vad som hände . 
Bara vinden och oljudet . 
- Det enda jag tänkte ... - Okej , Judy ... 
Det enda jag tänkte på var mina flickor ... Mina flickor skulle bli ensamma i världen . Utan mamma , utan pappa . Judy ! 
STREJKBRYTANDE BITCH 
Där är den . 
Hur känns den ? 
Vem skulle göra det ? 
Vem skulle göra det mot mig ? 
Gazza , någon ville döda mig , någon ville göra mina flickor föräldralösa . 
Hur kunde någon ... Hur kunde du ? 
Du . 
Du skar sönder mina däck . 
Du ville döda mig . 
HJÄRTAT BRISTER VI TÄNKER PÅ ER HÖGAKTNINGSFULLT , GAZZA MED FAMILJ 
Förlåt . 
Förlåt . 
Jag vill inte ha dina ursäkter . 
Vad fan tänkte du på ? 
Eller var det någon annan ? 
Gazza , du måste förklara , annars får du prata med polisen . 
Den skulle klara en bomb . 
Är du säker ? 
Vi har inte mycket tid . 
Jag går efter sovsäckarna , du går efter maten . 
Och sedan måste du göra dig klar för skolbalen . 
Jag tänker inte vara klädd som en jättelik maräng när världen går under . Okej ? 
Jag stannar här . - Gör det här rätt . 
- Du går på balen . 
Din mamma har sytt klänningen och Jono väntar på dig . 
Tilly , kom hit . 
Vi kan inte sluta leva . Fast vi är rädda . 
Du har aldrig varit så här rädd . 
Har du ? 
Nu säger de att Skylab kan störta här . 
Tilly och jag visste det redan . 
Lam , du oroar dig för mycket . 
För min familj , ja . 
" Tre omloppsvarv i dag . 
Den sista rakt ovanför Perth ... " 
Jag måste hålla dig säker . 
Det gör du . Lam , det har du alltid gjort . 
Skräm inte Binh , okej ? 
Det är hans och Tillys stora kväll . 
Jag meddelar markkontrollen . 
SISTA VARVET FÖR SKYLAB 
Jag har en överraskning till dig . 
Den är till din kostym till balen . 
Om Tilly är som pappa , kommer hon kanske inte . 
Jävla Skylab . 
HEMLIGSTÄMPLAD INFORMATION 
TILLHÖR KORPRAL GEORGE BARNES 
JAG SKULLE SKRIVA OM MIN DAG MEN JAG HAR GLÖMT DET MESTA 
NÅGRA KOMPISAR FICK LÄRA SIG OM FARORNA GÄLLANDE KÄRNVAPENTESTEN 
VI ANSER ALLA ATT DET ÄR SKITSNACK 
ANTHONY OCH GEORGE 
- Vi ses i kväll på balen , Rosie ! 
- Ja , vi ses där . 
Tony . Hur mår du ? 
Jag trodde du var upptagen med din kostym för i kväll . 
Tony ? 
I går kväll när jag hörde dig ... Din historia ... 
Jag visste inte att du var där . 
Jag beklagar . 
Jag var också där . 
Rekryterad . 
Jag ville glömma . 
Jag kan inte begrava det längre . 
Ville du glömma ? 
Jävla tur för dig . 
KVINNOR , INTE OBJEKT 
- Vad vill vi ha ? 
- Jämlikhet . 
- När vill vi ha det ? 
- Nu ! 
Fyra timmar kvar . Sedan kan de bränna bysthållaren och äta förbaskad falafel igen . 
VEM TILLHÖR DIN KROPP ? 
Hej . 
- Svetlana , det är jag . 
- Var är du ? 
Jag är på nedervåningen . 
Gäller det nu ? 
Ja , snart . 
Jag ringer när vi är redo . Då kommer du ner . 
Yvgeny kommer snart tillbaka från sin briefing . 
- Skynda . - Har du packat ? 
Har du allt du behöver ? 
Självklart har jag packat . 
Ring mig när jag ska komma . 
Var redo , hejdå . 
Det var snabbt . 
Nej . 
Han är inte här . 
Tack . 
Vad ? 
Vad är det ? 
Yvgeny , sätt dig . 
Vad är det ? 
- Har nyheten om babyn läckt ? 
- Nej . 
Om det bara vore det . 
Det var från Moskva . 
Din son ... 
Nikita ? 
I Afghanistan , hans grupp , den ... Hans trupp ... 
Jag är så ledsen . 
- För Guds skull , Jude , sluta oroa dig . 
- Jag oroar mig inte . 
Bara demonsonen inte står emot , är Murray hygglig . 
När han skötte affärerna var han rakt på sak . 
Allt ordnar sig . 
När det här är klart , är det vi som sköter affärerna , och vi lagar ett cocktailkabinett i Waynes gamla kontor . 
Varför är jag här ? 
Jag har ett företag att sköta . 
Du är en sakésvingande revolutionär , min vän . 
Fran ? Är du full ? 
På allvar . 
Eftersom Judy inte förstod sig på Japanska för nybörjare , är du för tillfället översättare . 
Du får visa hur Wayne urholkade företaget . 
Damer . 
Murray , detta är Hiroshi . Japansk översättare . 
Murray Doull . 
Hiroshi Hatano . 
Vad handlar det här om ? 
Dumme lille jävel ! 
Det är ett sätt att beskriva honom på . 
Johnnie Walker . 
Dubbel . 
Femtio år tog det att bygga detta företag . 
Men vi kan göra något åt saken . Vi måste göra något i kväll . 
Miss Universum och varningarna om Skylab , det är bara några timmar kvar , om det blir strömavbrott ikväll , och vi inte har löst dispyten , då är det kört för ditt företag . 
Det kommer inte finnas något att rädda , eller sälja . 
Vilket svek ! 
Att han skulle konspirera för att göra dig illa , Judy , för att få bra karlar att se dåliga ut . Att sätta dit facket , avskeda arbetarna och sälja oss utomlands . 
Flaskan . 
Detta japanska avtal , är det bindande ? 
Låter det honom sälja företaget utan arbetarna ? 
Det är i princip bara en överenskommelse . 
Okej , jag har klarat mig ur svårare lägen . 
Wayne får gå . Han klarar det inte . Jag är tillbaka . 
Fran , vi måste gå till facken . Nu ... Säg att det är från mig personligen . 
Släpp nyheten till pressen omedelbart . 
Jag tar hand om facken . 
Du måste ta hand om din familj . 
Du får gå . 
- Men chefen , jag tycker ... 
- Fran . 
Du får ett rejält avgångsvederlag , och min tacksamhet , men jag kan inte ha dig kvar efter att min son fått gå . 
Dags att gå vidare . 
Bob , knacka två gånger på fönstret om du ännu gillar mig . 
- Hej , mamma . 
- Åh , herregud . 
- Hur mår du ? 
- Jag är överraskad . 
Jag trodde inte vi skulle se dig på ett tag . 
Varför är du uppklädd ? 
Du ser jättefin ut . 
Jösses . 
Mamma ... 
Visst är han snygg ? 
Kolla vilken moodidj maman ! 
Är det så här du fostrar och stärker en ung man från ursprungsfolket , genom att klämma in honom i en jävla kostym ? 
Det är exakt därför jag kommit för att hämta min son , för att ta honom tillbaka till sitt folk . 
Jag ska gå på skolbalen med skolans häftigaste tjej , och hon valde mig för jag är den bästa dansaren . 
Mormor är mitt folk . 
Hon talade ut på radion , hon berättade för hela västra Australien , om oss och om morfar . 
Hon berättade sanningen . 
Alla hörde det , vi ... 
Vi har det på kassett . 
NANS SANNING 
Inlägget var så bra att de upprepade det . 
Lugna dig , mamma . 
Min kostym är inte som de andras . 
Vad fan händer ? 
Jag ringde dig som planerat , du skulle komma ner . 
Yvgeny ? 
Är han här ? 
Hans son var soldat i Afghanistan . 
Han dog för tre dagar sedan . 
Han är helt ensam , jag kan inte lämna honom . 
Det skulle krossa honom , det vore elakt . 
Jag har tjänstgjort . 
Jag förstår . Förlust . Men du är inte skyldig honom något . 
Bara dig själv . 
Kanske det är skillnaden mellan oss . 
Vi har våra brister . Men vi sätter inte oss själva först . 
Jag lämnar honom inte ensam . 
Han skulle inte göra det mot mig . 
Svetlana , om vi inte går nu kanske du inte får en andra chans . 
Han satt där , med ett whiskyglas i handen , och han sa , " Du ska ta hand om din familj . " 
Tio minuter , flickor . 
Kanske han borde gå och ta hand om sin avkomma . 
- Är det där ... 
- Min bröllopskostym , ja . 
Och ja , den passar än . 
Lite sliten , kanske . 
Den passar än . 
Liksom äktenskapet . 
Hur mår min familj ? 
Tilly kommer aldrig att jobba på jävla Boans . 
Hon tycks veta mer än NASA om Skylab . 
Och Mia försök hålla henne borta från surfandet . 
Och du ? 
Du vet hur jag är , hur vi alla är . 
Du behöver inte börja ta hand om din familj . 
Du har gjort det hela tiden . 
Men det visste du . 
Vad jag inte vet är vad som händer härnäst . 
Jag kan inte bara fortsätta . 
Jag kan inte gå tillbaka . 
Nej . Det ska du inte . 
Men jag måste gå tillbaka till Maralinga , jag måste berätta sanningen . 
Du ledde facket i 15 år . 
Du slogs för det goda , du din envise jävel . 
Du fixar det här . 
Ja . 
Och den där gamla saken ... 
Hallå ! Vet du vad fan din fru har gjort ? 
Jag har förlorat allt . 
Min pappa , mitt företag . Mina inkomster , tack vare din bitch . 
Nej , Tony . Tony , snälla . 
Var snäll och ta hand om flickorna . 
Jag sköter det där . 
- Du fattar inte , va ? 
- Upplys mig . 
Jag är inte bara Tonys fru . Och jag är definitivt inte hans bitch . 
Jag är ingens bitch . Och du är inte längre min chef . 
I själva verket är du ingens chef . Och den här tillhör dig . 
Du borde kanske be Gazza ge tillbaka dina pengar . 
Han visade sig vara en skitskytt . 
Gå bort från min gräsmatta . 
Och kom inte tillbaka , du din patetiske , lille pappas pojke . 
Fin kostym , pappa . 
Mycket stilig . 
Båda mina män . 
Stå tätt ihop . 
Perfekt . 
Okej . 
- Tre , två , ett . - Tre två , ett . 
Vänta tills jag berättar om hans kapten Stirling-byst . 
Gör plats åt pappa . 
Nu kör vi ! 
Se på dig . Du är en ung kvinna . 
Vad kvällen än betyder , njut av den . 
Okej ? Oroa dig inte för morgondagen , oroa dig inte för Skylab , oroa dig inte för något . 
Bara njut av kvällen . 
Skylab är i kväll . 
Den är antagligen ovanför Indiska oceanen just nu . 
Tilly . 
Tack , mamma . 
Och för klänningen , den är vacker . 
BITCH ÄR TILLBAKA 
Intrång ! 
Vi måste skydda våra flickor ! 
VI ÄR INTE OBJEKT SKÖNHETSTÄVLINGAR UTNYTTJAR KVINNOR 
- Vad vill vi ha ? 
- Jämlikhet ! 
- När vill vi ha det ? 
- Nu ! Sju minuter till ridå , flickor ! Sju minuter till ridå . 
- Släpp mig , släpp ! 
- Släpp mig . 
Klänningarna passar inte . 
Hela världen ser att jag är gravid . 
- Svetlana ... 
- Och i morgon , efter att jag kommer sist i kväll , är jag på enkel resa tillbaka till Sovjetunionen - och så är det med det . 
- Vi kan fly . 
Nu . 
Yvgeny klarar sig , det vet du . 
Vi ser efter varandra här . 
Jag har bevittnat det . 
På sätt som du inte kan tänka dig , i kriget , på gatorna , vi gör det . 
Stanna . 
Gift dig med mig . 
Se vad vi åstadkommit under de senaste veckorna . Tillsammans , inte ensamma . 
Vi kan göra det här , inte bara fly . Ett nytt liv . 
Det är garanterat bättre än att återvända . 
Sex minuter kvar , flickor ! 
Sex minuter . 
Jag kollar hur vi kommer härifrån . Jag är tillbaka om två minuter , okej ? 
Vad är det med honom ? 
Får jag presentera , Christine Baker . 
Den underbara Christine är i kväll tillsammans med Charlie , vicekapten i fotbollslaget Swan . Bra gjort , grabben ! 
Åh , den där klänningen . 
Stackars flicka . 
Det enda som är klumpigare än sömnaden är hans dans . 
Var försiktig , kompis , hon är en manslukerska . 
Till nästa , Mandy Barratts ... 
Tony ! 
Skylabs nästa varv börjar snart . 
Sista varv ? 
Ja , jag tror det . 
Varför är alla flickor klädda i likadana vita klänningar ? 
De ser ut som ledsna brudar . 
Vad ? 
De gör det ! Alla likadana . 
Se på dig . Du är inte likadan , va ? 
Okej . 
Du får surfa . 
Du ska surfa , men du måste också jobba , okej ? 
Du ska vara du . 
Det är allt . 
Ge en stor Scarborough-applåd till den vackra Becky Jones och hennes inhoppande partner , storebror Barry Jones ... 
Jones , vi tänker på dig och vi hoppas köttsåren läker snart . 
Vi älskar dig , Jones . 
Familjen som dansar ihop stannar ihop . 
Eileen . 
Vad vill du , Tony ? 
- Verkligen . 
- Eileen . 
- Jag menade inte ... 
- Ser jag ut som en präst ? 
Ber du mig om syndernas förlåtelse ? 
Eller vill du göra något åt det ? 
Den där skiten . 
- Det som hände där ute . 
- Jag måste göra något . 
Jag måste . 
Vi båda måste . 
Vi pratar . 
Ordentligt . 
Imorgon . 
Kom . 
Idag är Poppy i sällskap av den stilige Bilya Wilberforce . 
Vi ger dem en stor Scarborough-applåd ! 
Heja Poppy ! 
- Åh , nej ! 
- Du fångade henne fint , Bilya ! 
Charlie , här kan du få motstånd på fotbollsplanen . 
Charlotte Duffy ... allas favorit-engelsklärare . 
Det är en jävla skam . 
- Sluta . 
- Nej . 
- Sluta . Sluta . - Det vet du . 
Vad ? 
- Inget . 
- Pappa . Sätt dig . 
- Rocco , sätt dig . 
- Sätt dig , pappa . 
- Sätt dig . 
- Okej , Rose . Sätt dig ! Måste du ställa till en scen ? 
Vår skolas nätbollskapten Danielle MacDonald och hennes snygge kavaljer , Chris Shaw ... 
- Du ser fantastisk ut . 
- Tack . 
Är du nervös ? 
Nej , inte jag heller . 
Det är hela den här kvällen , det är ... löjligt . 
När som helst kan 70 ton smält rymdfarkost träffa oss ... 
- Tilly ... 
- Det är hela Perth . Borta . 
Och vi står här klädda som till bröllop . 
Jag borde vara i vårt skydd , tillsammans med min familj . 
- Har ni ett skydd ? 
- Ja , vi byggde ett . 
Knäppt , va ? 
Nej , inte alls . 
Min pappa har varit orolig hela dagen . 
Han lyssnar på nyheterna på radion . Kom , vi ser efter . Elaine Thompson är i kväll i sällskap av Jimmy Griffin . 
- Det måste ha hänt något . 
- Och till nästa Darlene White , som i kväll är tillsammans med den mycket stilige Steven Bates . 
Vi ger dem en applåd . 
Tilly har alltid varit ambitiös , men att gå på balen ensam - är kanske lite för mycket . - Det är Til . 
Tilly . 
Skylab kommer att träffa oss snart . 
- Jag sa att Skylab är på väg . 
- Gå bort från scenen nu . 
Jag kan inte längre klandras för det där . 
En rymdfarkost stor som ett höghus träffar oss inom en timme . 
Det är bara ett strömavbrott . Ingen anledning till panik . 
- Gå bort , nu . 
- För Guds skull . Jag ... Jag är nörden ni alla skrattade åt . 
Rymdnörden . 
Jag vet det här . 
Istället för att sitta här , borde ni söka skydd . 
Tilly har rätt . 
Skylab missade Indiska oceanen . 
Den kommer . Nu ! 
Ta skydd . 
Spring . 
Jag sticker . 
Damer och herrar , ingen panik . 
- Är det ett missförstånd ? 
- Det är vår flicka . 
- Håll er lugna . 
- Hon hade rätt . Lam . Kanske vi borde tömma salen . 
Gå in i bilen , vi går efter barnen . 
Vi har korsat oceanen , vi klarar det här . 
Binh ! Binh ! Du måste hitta Binh . 
Kom , vi måste ut härifrån . 
Gå , gå , gå ! 
Jono ! 
Vårt skydd , kom ! 
Jag måste göra något . På scen . 
Gå . 
Av alla rockstjärnor , varför han ? 
Bowie ? 
Kanske min vän inspirerade mig . 
Kanske jag är en Starman . 
Jono , Tilly . Kom . 
Gå . 
Två minuter till ridå , damer . Två minuter . 
Skylab . 
Darth Vader kan landa här i sina lårhöga boots , jag bryr mig inte . Showen fortsätter . 
Två minuter . 
Är du redo ? 
Jag är väldigt ledsen för din son , Yvgeny . 
Jag vet hur det är . 
Hur vet du det ? 
Nittio sekunder ! Nittio sekunder . 
Och jag är väldigt ledsen för det här . 
Väldigt ledsen , kompis . 
Spring ! 
Förlåt , Yvgeny . Jag kan inte gå tillbaka . 
Vad gör du ? 
Det är 45 sekunder till ridå . 
Vad gör du ? 
Pizza , Lydia . 
Vi ska gå ut och äta en jättelik pizza med en miljon kalorier ! 
Ditåt ! 
Du har 32 sekunder på dig att få flickan ut på scen ! 
Okej , vi klarade det . 
Mick . 
De är KGB . 
Det är bilen som följt oss . 
Nej , de är inte KGB . 
- Mick , de är KGB . 
- Lita på mig . 
Ni ASIO-killar är lätta att känna igen . 
Hon trodde ni var KGB . 
Men bara australier använder kortärmat på vintern . 
Jag heter Svetlana Natalya Kulkova och jag vill hoppa av till Australiska statsförbundet . 
Svetlana , snälla ! 
Stanna bilen ! 
Ni ASIO . 
Jag är Yvgeny Ilyich Pugo från KGB . 
Jag vill hoppa av . 
Vårt hemland har inget för mig längre . 
Nu kör vi ! 
Tack , miss Bermuda . 
Och nu miss Sovjetunionen ! 
Miss Sovjetunionen ! 
Jaha , vi går över till Donnie och den läckra miss Italien . 
Mamma , borde vi inte söka skydd ? 
Vet du vad , Djinda ? 
Jag är trött på att fly från saker som de vita ställer till med . 
Jag har fått nog . 
Vi är tillsammans . 
Vi tar det som det kommer . 
Pappa . 
- Kom . 
- Okej . 
- Har du hört från din bror ? - Självklart . Du ? 
Nej , och det vet du . 
Om berget inte kommer till mamma , måste kanske mamma gå och klippa till berget ? 
Gjorde du allt detta för mig ? 
Om jag kunde , skulle jag göra det . 
- Jag föredrog Toyotan . 
- Jag med . 
Jävla jänkarna . 
Vad är det egentligen du gör ? 
Jag ser efter henne . 
Jag ser efter honom . 
Jag gillar den här . 
- Kom ! 
- Tilly ! 
Mamma , pappa . 
Vad nu ? 
PRODUCENTERNA TACKAR RESPEKTFULLT ABORIGINERNA OCH FOLKET PÅ TORRES STRAIT-ÖARNA SOM ENLIGT TRADITION ÄGER MARKEN DÄR DETTA SPELATS IN , 
