Evigt ljus ? 
Evigt ljus ? Det är jag . 
Pike ... Nu om nånsin behöver jag dig . 
Pike Trickfoot . 
Jag har känt mig svag sen vi gick in i helvetet . 
Jag behöver veta att du ... Försoning existerar inte i de fördömdas rike . 
Avresans helveten är förbjudna . 
Men varför ? 
Om vi hittar Zerxus , får vi tag i reliken som vi behöver . 
Din själ är värdefull . 
Det finns de i helvetet som vill använda den för onda syften . 
Om du ignorerar mina ord lämnas du ensam . 
Vad betyder det ? 
Evigt ljus ? 
Vänta , snälla ! 
Pike ... Pike ? 
Pike ? 
Jag ropade ditt namn . 
Jag såg bara till att vi är omhändertagna . 
Skyddar din gudinna oss ? 
Ja . Absolut . 
Bra . För om vi ska klara det här , behöver vi alla sorters mirakel . 
Där är det , Hades stad . 
Okej . Hur ska vi göra ? 
Alla därnere är antingen demoner eller blir uppätna av en . 
Vi ser inte ut att höra hemma i helvetet . 
Såvida vi inte gjorde det . 
Lilleman ? Jaha . 
Dags att klä ut oss Dags att sminka oss Dags att bli jävligt läskiga - Ja , för fan . 
- Större horn . 
En kanin ? Kom igen . 
Okej , jag skojar bara , kompis . 
- Hur känns det ? 
- Grymt . 
Pike ? 
Kom . 
Är du okej ? 
Själarna . Jag önskar att jag kunde hjälpa dem . 
Keyleth hade kanske rätt . 
Är det värt att ta sig igenom helvetet för en relik ? 
Du hörde Raishan . 
Vi besegrar inte Thordak utan den . 
Allt med det här stället känns fel . 
Som att det är en synd att vara här . 
Vi kan nog inte vända . 
Det kommer att gå bra , kompis . 
Helvetet är inte så illa . 
Många har bett mig att dra hit . 
Vi måste gå . 
Scanlans förtrollning varar inte för evigt . 
Förlåt mig . 
Ni där . Ni ser inte bekanta ut . 
Vart ska ni ? 
Den fallna själen Zerxus Ilerez står i skuld till oss . 
Och vi vill inkassera den . 
Jaså ? 
Är ni modiga nog att träffa honom ? 
Vad fan ? 
Nåväl . 
Det var äckligt . 
Maten är klar . 
Vem står på tur ? 
Ni luktar annorlunda . 
Vi har inte badat på några tusen år . 
Ursäkta mig , vet ni var vi hittar Mässingsskallen ? 
Vi letar efter en som heter Zerxus . 
De var rädda för hans namn . 
Hitta mig . 
Vi går . 
Jag vill inte vara här längre än nödvändigt . 
Lag Draconia har det åtminstone lugnt i snön . 
Jag vidhåller att det hade varit säkrare att borra oss ut . 
Ja , men mitt sätt var coolare . 
Jag kunde gjort det coolt . 
Kima ! 
Hör du mig ? 
Kima ! 
Hon kan inte vara långt bort . 
Vad vill du göra ? 
Jag ska slita den jävla draken i bitar . 
Pike . Du ser för jävlig ut , även för att vara en demon . 
Jag tror att jag väntar här en stund . 
Ni kan fortsätta leta . 
Det är lugnt . Jag klarar mig . 
Sprid ut er . Men gå inte för långt . 
Jag gillar inte hur varelserna tittar på oss . 
All denna ondska . Evigt ljus hade kanske rätt . 
Vi borde inte vara här . 
Det är okej . Jag ska inte skada dig . 
Jag vill bara hjälpa dig . 
Befria den här kvinnan med ditt helande ljus . 
Pike ! 
- Vad händer ? 
- Min hjärna gör ont . 
Fan ! Scanlan , din förtrollning . 
Skriken stör min koncentration . 
Dödliga . 
Färskt blod . 
- Vi kan inte stanna här . 
- Du behöver inte upprepa det . 
Vi måste gå , Pikey . 
Skit . 
Var är den jävla Mässingsskallen ? 
Vi kan inte fly från en hel stad . Vi måste tillbaka till portalen . 
Inte utan skölden . 
De har blickar i skyn . 
Vad gör vi ? 
Den här vägen . 
Hörni , därnere . 
Ja ! Bra skådat , kompis . 
Var redo att hoppa ! 
Fan , det kommer att bli tajt ! 
Kliv in . 
Tack för hjälpen . Hoppas jag . 
Den här vägen . 
Vad är det här för ställe ? 
Snyggt trick . 
Vox Machina . 
Ni vet hur man gör en entré . 
Hur visste du att vi var på väg ? 
När man pratar om trollen ... 
Reglerna är unika i det här riket . 
Var försiktiga innan ni uttalar fler namn . 
Det var din närvaro jag kände . Varför sökte du upp mig ? 
Den riktiga frågan är : vad gör Evigt ljus präst här ? 
Vi skickades hit av J ' mon Sa Ord . 
Hen har lämnat nåt hos dig . Gryningsmartyrens sköld . 
Inte lämnat . Förlorat . 
Vad menar du med " förlorat " ? 
Varje årtionde kommer J ' mon för att testa sin dåliga tur vid mitt bord . 
Hen skulle inte ha satsat en sån artefakt , men rätt ska vara rätt . 
Jag antar att ni har nåt i utbyte . 
Ni kom inte till helvetet utan nåt annat än önsketänkande . 
Vad vill en djävulsman ha ? Guld ? 
För en relik ? 
Nej . Ni måste komma med ett exceptionellt erbjudande eller insats . 
Vill ni testa lyckan i spel ? 
Om vi vinner får vi skölden . Va ? 
Och om jag vinner , stannar du som min gäst . 
För evigt . 
Nej , Pike . 
Han kommer att fuska . 
Lugn . 
Regler är det som skiljer Avresan från existensens miserabla plan , likt ert . 
Fusk är inte tillåtet . 
Okej , vad är det för spel ? 
Vad i ... Pike ? 
Slå dig ner . 
Ett kontrakt ? 
För att se till att du inte får kalla fötter . Pike ! 
Nej ! - Är de ... 
- Trygga men tystade . Så att spelet förblir rättvist . 
Ska vi ? 
Så rent blod . 
Riktigt speciellt . 
Spelet heter Fem skallar . 
Varje spelare har fem kort , bestående av fyra röda och en svart skalle . 
När de har delats ut får du inte flytta dina kort eller röra motståndarens . 
Målet är att hitta min svarta skalle innan jag hittar din . 
Hur ? 
Varje omgång får man ställa en fråga som hjälp att hitta den . 
Men man måste svara sanningsenligt på alla frågor , annars får man ett hårt straff . 
Som jag sa , vi har regler här nere . 
Jäklar . De har schysta stolar i den här skithålan . 
Jag kan inte fatta att hon gör det . 
Om det är nån som kan genomskåda ett fulspel , så är det Pike . 
Det har sina fördelar att börja . 
Du är min gäst , så du får äran . 
Första frågan är din . 
Okej , då gallrar vi lite . 
Är din svarta skalle till höger eller vänster om ditt mittenkort ? 
Du känner inte Evigt ljus närvaro . 
Din frälsare är inte här , eller hur ? 
Det var inte min fråga . 
Till höger . 
Längst ut , det är ditt kort . 
Tyvärr inte . 
Men jag lärde mig nog mer än vad du gjorde . 
Alla har nåt som avslöjar dem om man gräver djupt nog . 
Ska du inte fråga mig nåt ? 
Dina vänner förlitar sig på dig . 
Du måste vara stolt över att alltid rädda dem . 
Det är inget kortspel . Han visste exakt vem han ville spela med . 
Jag försöker förstå reglerna . 
Säg mig , du heliga . Fick du ett val ? 
En väg att gå ? Va ? 
- Vi väljer inte ... - Vi väljer inte ... 
- Alla kan vara heliga . - Alla vägar kan vara heliga så länge man går den sanningsenligt . 
Ja , jag fick ett val . 
Fast valet var en lögn . 
Båda vägarna ledde till samma slut . 
Jag gavs ett liknande val en gång . 
Det kostade mig min familj . 
Min gud förrådde mig . Och det kommer din med att göra . 
Nej . 
Du försöker ta dig in i mitt huvud . 
Det kommer inte att gå . 
Jag har redan det jag behöver . 
Du har redan avslöjat dig . Dina ögon . 
Ditt svarta kort ? Andra kortet från ditt vänster . 
- Nej . 
- Kompis ! 
Det här är skitsnack . 
Du ändrar ämne . Du fuskar ! 
Hur ? 
Alla svar var sanningsenliga . 
Kontrakt eller inte , det här är en fars . 
Minikuken har rätt . 
Jag tänker inte se på längre ! 
Vänta , du kanske inte ska ... Dumma bekväma stol ! 
Pike Trickfoot , du är nu bunden till den här helgedomen i den Fallna riddarens tjänst ... i evighet . 
Vänta ... 
Snälla , du måste ge mig en chans till . 
Vad mer har du att erbjuda ? 
Va ? 
Det kan hon inte . 
En meningsfull insats . 
Fast jag har tyvärr ingen användning av den . 
För Gryningsmartyrens sköld behöver jag nåt mer betydande . 
Dina vänners själar . 
Nej , inte dem . Jag kan inte . 
Är din tro inte stark nog ? 
Okej . 
En omgång , vinnaren får allt . 
Vänta . Är vi insatsen ? 
Det känns så . 
Pikey ? 
Jag förstår varför Evigt ljus gynnar dig . 
Du är lika vårdslös mot dina nära som mot dig själv . 
Men den här gången börjar jag . 
Min tur . Min fråga . 
Det är nåt annorlunda med dig , Pike . 
Du är speciell . 
Har du nånsin undrat om Evigt ljus behöver dig mer än du behöver henne ? 
Det har aldrig slagit mig . 
Två kort ? 
Ljuger för dig själv . 
Oj , det var nytt . 
Det är inte rättvist . 
Sanningen är sällan det . 
Du har gjort det enklare för mig . 
Visa kortet till mitt höger . 
Synd . Din tur . 
Okej . Lägg ner skitsnacket . 
Vilket kort är din svarta skalle ? 
Intressant taktik . 
Jag säger det eftersom jag inte kan ljuga . 
Det är det i min hand . 
Längst till vänster . 
Två kort . 
Vad ska jag fråga nu ? 
Jag vet . 
Undrar du nånsin om ditt liv vore bättre utan Evigt ljus ? 
Ja . 
Det låter inte lojalt . 
Ditt vänstra kort . 
Spelet verkar nästan vara över . 
Skit . 
Gör mig en tjänst innan du vinner . 
Om du håller kvar mig här för evigt , förtjänar jag att få veta vem du är , vem du var och varför du valde mig . 
Okej . 
Se det som en sista eftergivenhet . 
Jag kommer från en tid för tusen år sen ... Då gudar vandrade bland de dödliga och värden styrdes av magi . Jag , som du , skyddade mitt hem som Första riddare . 
Medlem i Mässingsringen , en grupp som liknande din . 
Och precis som du trodde jag det bästa om dem . 
Jag var förblindad då mina vänner fördömde vår civilisation med sin nyfikenhet och hybris . 
Menar du katastrofen ? 
Gudarna startade krig mot Exandria . Och i kaoset mötte jag Plågans herre själv . 
Men han gav mig ett val istället för att döda mig . 
Dö med de andra , eller ansluta mig till honom och skona min familj . 
Jag trodde att om jag hade nog med tid , skulle jag kunna nå honom , rädda honom , tämja hans våldsamma hjärta . 
På grund av min dårskap , såg jag min man och son blekna med tidens påfrestningar och tappa alla minnen av mig . 
Som om jag aldrig hade existerat . 
Litade du på en bedragar-gud ? 
Självklart . 
Precis som du enfaldigt litar på Evigt ljus . 
Men det är ingen skillnad på gudar där ovan eller nere . 
Alla ljuger ! 
Jag beklagar alla du har förlorat . Men mina vänner är inte så och inte min gud heller . 
Ge det tid . 
Nu har vi ett spel att avsluta . Och du har en fråga att ställa . 
Okej . Jag tror att jag har det . 
Önskar du att din familj var här ? 
Va ? 
Du valde det här livet för att skona din man och son . 
Du säger att du älskade dem , men jag hör bara ånger . 
Så vill du ha dem hos dig i den här mardrömmen ? 
Eller är det för själviskt ? 
Jag ... Svara på min fråga . 
Önskar du att de var här och led med dig ? 
Nej , jag ... - Svara mig ! 
- Självklart inte ! 
Jag vet inte ens om du vet att du ljög . 
Nej . 
Och nu är mitt val mycket lättare . 
Som sagt , alla har nåt som avslöjar dem om man gräver djupt nog . 
Det kortet . 
Snyggt spelat , Pike Trickfoot . 
Det var lömskare än jag förväntade mig . 
Vi har alla blinda fläckar . Även du . 
Det är ovanligt att jag förlorar i min domän . Men jag accepterar förlusten . 
Ja , kompis ! 
Ja ! Se på det . 
Tacka gudarna . 
Jag antar att Evigt ljus ställde upp . 
Ja . 
Får bara Pike en souvenir ? 
Jag glömmer inte din historia . 
Tack för att du var en god förlorare . 
Jag glömmer inte din . 
Okej . Är nån annan redo att dra härifrån ? 
Definitivt . 
Här , ta det här . 
Det har mitt märke . Ni behöver det för att ta er ut säkert . 
Yenk , visa dem till dörren . 
Och hälsa så gott till J ' mon . 
Jösses , det var nära ögat . Hon har ingen aning om vad som flyter genom hennes vener . 
Det kvittar . Ett frö av tvivel har såtts och det kommer att fylla henne med hämnd medan vi ser det växa . 
Dina order ? 
Låt henne vara . Döda resten . 
Vi är hans släktingar . 
Tiden för hans uppstigning närmar sig . 
Det blir mycket lättare att ta sig ut än in . 
Bra . För jag kan inte äta fler kryp . 
Vad är oddsen att det inte är menat för oss ? 
Jag säger 50-30 . 
Vox Machina ! 
Jag hatar matte . 
