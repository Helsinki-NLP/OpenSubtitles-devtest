Det är vad alla kallar mig , som ett tecken på kärlek och respekt . 
Samsik eller farbror Samsik . 
Jag älskar det . Jag älskar mitt smeknamn . 
Kapitalförsvarsenhetens hemliga bunker 
Vi har några frågor . Det går fort om du samarbetar . 
Trevligt att se dig överste . 
Hanmin . 
San , är det du ? 
Är du också här ? 
San ! San ! 
Vi planerade inte det här ! 
Det var Samsiks fel ! 
Kan du prata med dem ? 
Säg att det var Samsiks fel ! 
Känner du till Sail Utvecklings vd Pak Doochill ? 
Ja . 
Du kallade honom Samsik ? 
Ja . 
Vad betyder det namnet ? 
Att hans folk fick tre måltider även under kriget . 
Vare sig det var hans familj , vänner eller släktingar lät han ingen gå hungrig . 
Uncle Samsik 
Uncle Samsik 
Tre måltider om dagen 
26 november 1959 Seoul , Sydkorea 
Amerikanska arméns oljeförråd 
- Två ? 
- Två . - Tjugotusen hwan . - För oljan . 
Vad heter " olja " på engelska ? 
Det är tio sedlar . 
Olja . 
Det är 20 000 hwan . 
Det är 20 000 hwan . 
- Lite till . 
- Vad fan säger han ? 
- Stick härifrån ! 
- Spring ! 
Vad hände ? 
Gu Haejun och Han Soo Seodaemunligan 
Fan . 
30 november 1959 Seoul , Sydkorea 
Rhee Seungmin ställer upp i omval 
Vi måste skydda president Rhee ! 
Samsik har kontakter överallt . 
När Gunsankillarna åkte fast för smuggling - fick Samsik ut dem . 
- Du har sagt det . 
Har jag ? 
Käftar du emot , din usling ? 
Våra killar skickades till Counter Intelligence Corps . 
Hur länge måste vi vänta ? 
- Tyst . - Jösses . 
Ni kan gå in nu . 
President Rhee är vårt hopp ! 
- Vårt hopp ! - Vårt hopp ! 
Ställ upp i omvalet ! 
- Ställ upp ! - Ställ upp ! 
Hej , kom in . 
Ställ upp i omvalet ! 
Farbror Samsik ? 
Vi stöder president Rhees omval ! 
- Vi stöttar ! - Vi stöttar ! 
Kom in . 
- Är ni med Seodaemunligan ? 
- Ja . Ni stal olja från USA:s armé . 
Ja , våra killar skickades till CIC . 
Varför CIC ? 
Ingen aning . 
I Osaka äger ligamedlemmar bilar . Så hur kommer det sig att ni bara snattar ? 
Gör nåt med lite mer substans , okej ? 
Berätta . Kan du få ut våra killar eller inte ? 
Vad får jag ut av det ? 
Vi belönar dig rejält . 
Du är rätt kaxig för nån som ber om en tjänst . 
Vi drar . 
Var inte sån , Han Soo . 
- Vi går . 
- Så gulligt . 
Ska du bara gå ? 
Testa att kalla mig farbror Samsik . 
Pratar du med mig ? 
Kalla mig farbror Samsik . 
Varför skulle jag ? 
Då ger jag dig mat . 
Det gör dig inte till min farbror . 
Du vet Yoon Palbong från Dongdaemunligan ? 
Vill du ha hans område ? 
Han är med liberala partiet . Så hur kan vi ... 
Jag ger er det . 
- Fröken Kim , ge mig tio kuvert . - Ja ? 
Ta pengarna och bryt Yoon Palbongs ben . 
Protester mot president Rhees avhopp fortsätter över hela landet . 
Politiska kretsar övervakar noga om president Rhee kommer att svara på folkets begäran - och ställa upp för omval . 
- Kom , Jina . 
Jina . 
- Vi måste skydda president Rhee ! Farbror San , blir vi rika om det här utförs ? 
Studera hårt , okej ? 
Ta på dig skorna . 
Vi går nu . 
- Ha en bra dag . 
- Kom . 
- Vi ses , Jina . - Vi ses , mamma . 
Inrikesministeriet 
Rekonstruktionsbyrån . Hej , hur är det ? 
Herr Kim . 
- Ja ? - Telefon till dig . 
Vem är det ? 
Kim San från Rekonstruktionsbyrån . 
- Hej , San . 
- Yeojin . 
Passar det nu ? 
Ja , varsågod . 
Du borde inte komma i dag . 
- Det har snokats på sistone . 
- Snokats ? 
Jag kommer efter jobbet . Oroa dig inte . 
Vi ses sen . 
Herr Kim , ministern kommer . Skynda dig . 
- Ja , herrn . 
- Fröken Kim . 
- Ja ? Seohae oljas fabriksområde 
Ser du Seohaes oljefabrik från där du är ? 
Ja . 
När den är byggd blir jag officiell medlem i Cheongwooförbundet . 
Vet du vad det betyder ? 
Du blir den koreanska adeln ? 
Adeln , knappast . 
Jag blir den som störtar adeln . 
Kom igen . Skynda . 
Kom igen . 
- Han kommer nu . Skynda . - Okej . 
General Jang möter dig vid Taepyeonggak . 
Vad ska han proppa i sig den här gången ? 
Bra jobbat med skorna . 
Här kommer Yoon Palbong . 
- Fortsätt gå . 
- Hallå , Samsik ! Ignorera honom . 
Vänta , Samsik ! 
Herregud . Hur mår du , herr Yoon ? 
Jag samlar ihop 25 killar sen . 
Det känns verkligen betryggande . 
Pratade du med Kang Seongmin ? Det gjorde jag . 
- Du . 
- Kom igen , folk tittar . 
- Prata ordentligt . 
- Ställ inte till med en scen . Om det vi gjorde i Busan kommer ut är vi och Kang Seongmin döda . 
Han måste få mig nominerad för Dongdaemun . 
Är du galen ? 
Bad jag dig inte hålla tyst om Busan ? 
Jo , om Kang Seongmin håller sitt löfte . 
Varför är du så otålig ? 
Ledamot Kang har planerat allt . 
Varför undviker han mig ? 
För att du är överallt . 
Tänk på vad vi gjorde för honom . Men vi fick inget tillbaka . 
Jag ska visa vem som bestämmer på Innovationspartiets tal . 
Säg att det här är hans sista varning . 
Den jäveln måste vara galen . 
Avlägsnade du poliserna ? 
Ja , jag ordnade det . 
Idioten kommer att göra bort sig . 
Då sätter vi igång . 
Arbetslösheten skjuter i höjden på grund av kollapsen av småföretag , tillverkare och bönder . 
Jordbruksöverskott från USA driver på jordbruksskulderna . 
Med 80 % av skulden i privatlån med 6 % ränta , är jordbruksekonomin nära kollaps . 
Med vår unga arbetskraft ... 
Presidenten frågar efter dig . 
Ställer han upp i valet ? 
Det är inte säkert än . 
- Det var allt . 
- Genomgången har bara börjat . 
- Vi ses . 
- Mitt team jobbade hela natten . 
Vem är han ? 
Rekonstruktionsbyråns chef , Kim San . 
Herrn . 
Koreas framtid ligger här . 
Vem tror han att han är ? 
Han studerade ekonomi i USA med ett Albrightstipendium . 
- Albright ? - Ja , herrn . 
- Gick du på militärakademin ? 
Vad gör du här ? 
Passade du inte i armén ? 
Herrn , presidenten väntar . 
Skicka en rapport . 
Jag har skickat flera . 
Vi skickar den igen . 
Jag har gjort det i två år . 
Presidentvalet är vår högsta prioritet nu . 
Vem bryr sig om det ? 
Arbetslösheten är hög , jordbruksekonomin är död , och vi behöver USA:s stöd . 
Är han galen eller ? 
Ge mig en timme , herrn . 
Herrn . 
Herrn ! 
Bara en timme ! 
Herregud . 
Vi har skickat rapporter i två år . 
Taepyeonggak 
- Sjöfågel - Sjöfågel 
- Varför gråter du ? - Varför gråter du ? 
- Förakta inte tiden - Förakta inte tiden - Som flyger förbi ... - Som flyger förbi ... 
Sjöfågel 
Varför tog han med så många ? 
Ingen aning . 
- Livet går och kommer ej åter - Livet går och kommer ej åter - Kvar blir de gröna bergen - Kvar blir de gröna bergen 
Du , Samsik . 
Märkligt . Vart tog spriten vägen ? 
Det var hit upp . 
Vad gör en general här med nybörjarna ? 
Man kan inte vinna deras lojalitet utan att bjuda dem ibland . 
Men det är jag som betalar . 
Känner du Hong Youngki , chefen för CIC ? 
Hong Youngki ? 
Varför ? 
Min brorson sitter på CIC för att ha stulit olja från USA:s armé . 
Vill du få killarna släppta ? 
Nåt i den stilen . 
Är det nåt man ber en general om ? 
Det var därför jag gjorde dig till general . 
Vet du inte hur Hong Youngki är ? 
Inte ens en general kan göra mycket under hans uppsikt . 
Förra året sparkade han en tredjedel av generalerna . 
Hur ? 
Han kan märka vem som helst som kommunist . 
Han kokar ihop bevis och burar in dem . 
- Han låter som jag . - Vad menar du ? 
Om han kan sparka en tredjedel av generalerna , varför skulle han bry sig om småtjuvar ? 
- Han använder dem som lockbete . 
- Lockbete ? 
Prata med honom . 
Är du galen ? 
Gå emot ministern ? Varför inte slå honom i ansiktet ? 
Om du vill få som du vill , ge dig in i politiken ! 
Gå i herr Choo Intaes fotspår ! 
Kampanja , håll tal , eller vad som helst ! 
- Det ska jag . 
- Va ? Jag ska hålla tal om aktuella frågor sen . 
En statsanställd som håller tal på Innovationspartiet ? 
Herr Choo är som en far för mig . 
- Han är inte din riktiga far ! 
- Jag går nu . Hallå ! 
Du kan inte gå under arbetstid . 
Jag är trött på rapporter . 
Skriv den inte . 
Presidentens kontor 
Det är min tredje mandatperiod som president . 
Det är folkets önskan . 
Jag drog tillbaka min kandidatur . 
Folk skulle håna mig ... " President " ... om jag gör tvärtom . 
Har du sett Choo Intaes popularitetssiffror ? 
Har jag en chans mot honom ? 
Jag gör vad som helst för att du ska vinna . 
Vad som helst ? 
Ja . 
Du kan vara lugn . 
Hotell Banya 
Efter vägledning från Cheongwooförbundets medlemmar ... 
Ja , hej . 
Nu ska vi se . Fortsätt så . 
Efter vägledning från Cheongwooförbundets medlemmar har jag äran att stå här i dag . 
" Har jag äran ... " Så töntigt . 
Så ? 
Är du redo ? 
Jag är så nervös . 
Grattis . 
Alla får inte gå med i Cheongwooförbundet . 
Det betyder att du är en av landets 20 bästa affärsmän . 
Tack vare herr An Yosubs vägledning har jag äran att stå här i dag . 
När vårt industrikomplex är klart får vi äntligen äta pizza som amerikanerna . 
Ni har nog aldrig hört talas om pizza . 
Det är jättegott . 
Nog med prat . 
Genom att säkra en andel på 60 % i Seohae Olja , får nu Samsik ... jag menar Pak Doochill , 
Accepterar vi honom som ny medlem ? 
Petron Harvest , Sierra Union , Hassel Chemistry ... 
Alla åtta potentiella partners gav samma svar . 
De kräver betalningsgarantier från regeringen , rätten att använda hamnar , kontroll över järnvägen och diplomatstatus för industrianställda ? 
De kan avbryta affären ! 
An Kichul An Yosubs yngste son 
Vet du vad pizza är ? 
Det gör du säkert inte . 
Ugnen är större än ditt sovrum och brödet är lika stort som du . 
Det toppas med kött , ost och grönsaker . 
En tugga och ... 
Du vet nog inte vad ost är heller , va ? 
Ost ? Nåt slags bröd ? Jösses , så typiskt för en kroppsarbetare . 
Du vet ingenting , va ? Hur lyckades du gå med i Cheongwooförbundet ? 
Amerikaner äter sånt bröd varje dag . 
Ibland äter de inte upp . 
När vårt industrikomplex är klart blir vi både mätta och kan slänga lite . 
Det måste finnas en anledning till att de gör så . Tänk på vår investering i industrikomplexet . 
Det är konstigt att alla åtta gör det samtidigt . 
Jag ska ta reda på deras avsikter . 
Kang Seongmin . 
Jag vill ha hit honom nu . 
Ja , herrn . 
Den dagen kommer . 
Hur gick det ? 
Vad är det ? 
Petron Harvest har fler krav . Va ? Vad för krav ? 
Det är på engelska . Jag kan inte läsa . 
De vill ha betalningsgarantier från regeringen , rätten att använda hamnar och övervaka statliga bidrag . 
Var kommer det här ifrån ? 
De kan nog inte lita på vår regering . 
Vad händer nu ? 
Vad tror du ? Våra planer kan gå i stöpet . 
Jag då ? 
Jag gick precis med i förbundet . 
Det går inte utan Seohae Olja . 
Hördu , ut med dig . 
Ledamot Kang . 
Varför är det så svårt att nå dig ? 
Jag bad dig sluta dyka upp . 
Hörde du om Innovationspartiets tal ? 
Jag skickade 25 killar till . 
Äras den som äras bör . 
Visst . 
Vi pratar efter presidentvalet . 
Ryktet säger att nån annan kommer nomineras till Dongdaemun . 
Sluta utnyttja mig och håll din del av avtalet . 
An Yosub är väl därinne ? 
Ska jag berätta vem som dödade hans son ? Tänk om han får veta vem som dödade An Minchul i Busan . Vad tror du han gör då ? 
Kang Seongmin Liberala partiets ledamot 
Det här har varit vårt mål hela tiden . 
Om industrikomplexet misslyckas behöver vi en plan B. 
Du är här . 
Kan vi prata , farbror Samsik ? 
Jösses . Du verkar bekymrad . 
Yoon Palbong besökte mig igen . 
Va ? 
Igen ? 
Jag pratade ju förstånd med honom . 
Jag ska lära honom en läxa på Innovationspartiets tal . 
Oroa dig inte . 
Döda honom . 
Ursäkta ? 
Döda Yoon Palbong . 
Så fort som möjligt . 
Jag är livrädd . 
Jag drömmer om den döde An Minchul . 
Yoon Palbongs högsta önskan är att bli ledamot . 
Kan han inte få bli det ? 
Döda honom bara . Jag kan inte fortsätta så här . 
Okej . 
Som du vill . 
Du är allt jag har , farbror Samsik . 
Hjälp mig att sova på natten . 
Alla åtta potentiella partners skickade in de här . 
Varför nu ? 
De tycker att vår regering är opålitlig . 
Varför tror du att jag gjorde dig till ledamot ? 
Om Minchul fortfarande levde , skulle han sitta där du sitter nu . Han hade gjort ett bättre jobb än du . 
Kang Seongmin vill att jag dödar Yoon Palbong . 
Varför ? 
Yoon Palbong pratar om Busan hela tiden . Om hur vi dödade An Yosubs son . 
Tror du presidenten ställer upp för omval ? 
- Inget är säkert ... 
- Det gör han . 
Han anlitade till och med demonstranter . 
Jag kollar upp det . 
Du är alltid ett steg efter . 
Våra planer för industrikomplexet kan gå i stöpet . 
Kang Seongmin är en fegis . 
Han kan inte slappna av förrän allt och alla han är rädd för är borta . 
Menar han allvar om Yoon Palbong ? 
Jag blir hans nästa mål . 
De med makt och pengar smutsar aldrig ner sig . 
Varför tror du att han bad mig döda Yoon Palbong ? 
Jag har känt Kang Seongmin sen han var liten . 
Han har en speciell min . En elak , kallhjärtad min . 
Hans min när han bad oss döda An Minchul . 
Han hade samma min nu . 
Vänta och se . 
Han försöker säkert döda mig härnäst . 
Petron Harvest skickade ett inspektionsteam till Filippinerna . 
Planerar de att utföra våra planer där ? 
Det är möjligt , med tanke på inspektionsteamet . 
Vi gör allt jobb och nån annan får äran . 
Choi Minkyu tog för lång tid på sig . 
Jag pratar med ministern . 
Säg att vi är redo att möta alla krav . 
Yeojin . 
San , du är tidig . 
Hur går förberedelserna ? 
Jag gör mitt bästa , men jag är osäker . 
Min far har aldrig talat till allmänheten . 
Oroa dig inte . 
Det går nog bra . 
Hitåt , minister Choi . 
Seonyoowon 
Minister Choi är här . 
Han är framme i Seonyoowon . 
Yoon Palbong skickar 25 män till Innovationspartiets tal . För att föra liv under herr Choo Intaes tal . 
Han har gjort det under det senaste årtiondet . 
Han har attackerat oppositionspolitiker på nåns order . 
Hur stort är ditt gäng ? 
Vi är 15 personer . 
Klarar ni av 25 personer ? 
Haejun , Heesung och jag är i korridoren . 
Jongsol , omringa Dongdaemunkillarna med lastbilen . Mer chilipulver . 
Att ta sig an 25 personer är enkelt , men efteråt , då ? 
Polisen griper bara oss och inte Dongdaemunkillarna . 
Om jag avlägsnar poliserna , då ? 
Kan du göra det ? 
Undan . 
Är det inte uppenbart ? 
Han Soo , polisen drar sig undan . 
- Allihop ? 
- Ja . 
I så fall kan vi lätt ta oss an 25 personer . 
Yoon Palbong får inte komma undan . 
Se till att bryta hans ben , okej ? 
Det blir en folksamling vid Choo Intaes tal . 
Förutom ledamöter , kommer alla möjliga att vara där för att smöra för Choo Intae . 
Han är populärare än presidenten just nu och kommer nog att vinna valet . 
Därför är han en måltavla . 
Choo Intae Innovationspartiets ledare 
Innovationspartiets tal 
Fredlig återförening och vår nations väg av Choo Intae 
Jag vill välkomna alla till Innovationspartiets tal om aktuella frågor . 
- Choo Intae ! - Choo Intae ! - Choo Intae ! - Choo Intae ! 
Tack , allihop . 
Jag är Choo Intae . 
Vilken väg ska nationen ta ? 
Vår prioritet borde först och främst vara en fredlig återförening och samexistens mellan Nordkorea och Sydkorea . 
- Ja ! - Ja ! 
Vad har den nuvarande regeringen gjort för folket hittills ? 
Absolut ingenting förutom att ödelägga böndernas och arbetarnas liv . 
- Ja ! - Ja ! 
Hördu . 
In med dig , för fan . 
Fan , lycka till . 
Den sittande presidenten visar upp sig genom att dra tillbaka sin kandidatur . 
Vem går på det ? 
Ja ! - Ja ! - Ja ! 
Det är flera Dongdaemunkillar i korridoren . 
Kan du ta dig an dem ensam ? 
Självklart . Bara säg var de är , farbror Samsik . 
Hur kan han sjunka så lågt ... 
Kör . 
... för att bli omvald ? 
Han insisterar på återförening genom att störta Nordkorea ! 
Men vem betalar priset för det ? 
Tänk er 100 män var . 
Minst tre män var ! 
Det här landet ska aldrig behöva uppleva ett krig igen ! 
- Choo Intae ! - Choo Intae ! - Choo Intae ! - Choo Intae ! 
Choo Intae är kommunist ! 
Hallå ! 
Era jävlar ! 
Följ med mig . 
Ring polisen ! Skynda ! 
- Hallå ! - Vem är du ? 
Ring polisen . 
Ring den jävla polisen , sa jag . 
Kom ut när du har skitit klart , idiot . 
Jag gjorde det , eller hur ? 
Nu drar vi . 
Förresten , har herr Choo redan rymt ? 
Kan en så feg kommunist hantera politik ? 
Precis . 
Ursäkta mig . 
- Pratar du med mig ? 
- Vem är du ? 
Ledamot Pak från Liberala partiet . Du borde sluta . 
Lugna dig , ledamot Pak . 
Lugna dig . 
Vem är du att tilltala en ledamot så ? 
Herr Choo är inte kommunist . 
- Be om ursäkt nu . - Va ? 
Herr Choo står för nationens välstånd och fredliga samexistens . 
Det låter precis som en kommunist . 
Vet du hur han är ? 
Har du läst Framgång på Koreahalvön ? 
Den utforskar vårt folks ekonomiska pånyttfödelse . 
Det visste du nog inte . 
- Nej . Idiot . - I så fall , får jag förklara det ? 
- Varsågod . 
- Tack , herrn . 
Låt oss lyssna . 
Jag kommer hit när jag känner för att ta en drink ensam . 
Kom gärna hit och ta en drink när du vill . 
Handlar det om industrikomplexet ? 
Det är hopplöst . 
Presidenten är emot det . 
Enligt honom är planerad ekonomi kommunistiskt . 
Hej , allihop . 
Jag jobbar på Rekonstruktionsbyrån . Jag doktorerade i ekonomi i USA . 
Jag har varit i USA som Albrightstipendiat . 
I USA var allt överflödigt och vackert . Men mitt land var slitet och mitt folk svalt . 
Vet nån vad pizza är ? 
Har nån smakat det ? 
Har du smakat det ? 
Nej , din lilla snorunge . 
Jag bodde ovanför en pizzeria i USA . Jag åt knappt en måltid om dagen . 
Doften av pizza höll mig vaken om natten . 
Ekonomin kommer före vapen och svärd . 
Ett land där ingen går hungrig och där alla kan få tre måltider varje dag . 
Det jag avundades mest i USA var varken stridsflygplan eller hangarfartyg . Det var pizza . 
Varför vinna ett krig om alla i landet svälter ? 
Det var då herr Choo föreslog att jag skulle studera ekonomi . 
Stål , skeppsbygge , transport , kemikalier , olja och textilier . 
Alla landets nyckelindustrier . 
Cheongwooförbundets medlemmar har satsat allt på detta . 
Om vi missar denna chans förlorar vi alla våra partners till Filippinerna eller Taiwan . 
Vi kan inte investera mer i anläggningarna . 
Vi har redan lagt alla våra pengar på dem . 
Utan utländskt kapital är våra investeringar förgäves . 
Så om regeringen kan hjälpa oss ... 
Vad händer då ? 
Ska du hjälpa oss i presidentvalet ? 
Ja . 
Både presidenten och herr An Yosub är över 80 . 
Hur länge tror du att de sitter kvar vid makten ? 
Jag står på tur . 
Efter mig kan det bli du . 
Din förmögenhet och bakgrund och min makt . 
Vad tror du händer om vi delar det vi har ? 
Jag tror att vi blir oövervinnliga . 
Visst , jag antar det . 
Använd presidentvalet för att ta kontroll över partiet . 
Bli valkampanjens ordförande . 
Det är klart när jag frågar presidenten . 
Jag ger dig chansen att ta kontroll över Liberala partiet . 
I så fall vad ska jag ge dig i gengäld ? 
Cheongwooförbundet . Vad annars ? 
Titta på det här . 
Vi ska bygga en motorväg mellan Seoul och Busan , upprätta industrikomplex och hamnar , bygga en motorväg mellan Seoul och Incheon och exportera varor från Incheon till Kina . 
Kina har 700 miljoner invånare . Om varje person köper ett par skor säljer vi 1,4 miljarder skor . 
Din idiot . 
Varför skulle vi sälja skor ? 
Du låter som en kommunist . 
- Ja ! - Ja ! 
Har inte kommunister skor ? 
Just nu med vår unga arbetskraft , kan vi bli en industrialiserad nation . 
Med tre hav inom räckhåll kan vi få ett övertag i handeln . 
Det är det landet herr Choo drömmer om . 
- Choo Intae ! - Choo Intae ! - Choo Intae ! - Choo Intae ! 
