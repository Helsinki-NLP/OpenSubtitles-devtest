Nej ! 
Återgäldar ni mitt överseende genom att attackera min tron ? 
Jag ska förvandla er till aska . 
Få bort männen härifrån . 
Det här är illa . 
De kom för att hjälpa oss och nu ... De blir slaktade . 
Thordak skulle inte lämna sina ägg . 
Vi skulle överraska honom . 
Herregud ! 
Vi kan inte stanna här , vi måste göra något . 
Det finns inget vi kan göra . 
Där sket sig den planen . 
Har någon en annan plan ? 
Percy hade haft en plan . 
Resten av äggen kläcks snart . 
Jag tycker vi följer strategin . Tar oss till nästet medan armén är vid fronten . 
De skulle bara slåss mot de små , inte Thordak ! 
Och Raishans tunnel finns inte . 
Vi tar oss inte in . 
Vi har huvudingången . 
Den som Thordaks barn vaktar ? 
Den som vi sa var för farlig ? 
Vi kan inte lämna de andra . 
Thordak dödar dem på två minuter . 
Vår hjälp kan förlänga det med en minut . 
Åt helvete med det här ! 
Vi gör båda delarna . 
Keyleth , Pikey , hjälp armén . 
Tvillingarna ansluter när jag och Scan är i nästet . 
Vi krossar äggen , ni krossar hans kristall . 
Några frågor ? 
Det var imponerande . 
Förlåt , jag fick en blackout . 
Vad sa jag ? 
Kom igen , snillet , nu flyger vi . 
Ballister , skjut ! 
Gör ditt bästa , byracka . 
Fri eldgivning . 
Jag har dig . 
Vad hände ? 
Vad gör ni här ? 
Vi ville inte att ni skulle dö ensamma . 
Det är ... Det är ett dåligt skämt . 
Vi måste få bort soldaterna härifrån nu ! 
Vart då ? 
Vi ger oss på Thordak och håller honom sysselsatt . 
Du fördömer oss . 
Vi borde ta oss an de små för att ta oss fram . 
Fattar ni inte ? 
Vi är instängda utan utväg . 
Vad sa du , vännen ? 
Genom den väggen , fort . 
Kom ! Zahra ! 
Kash ! 
Ni skulle inte komma . 
Jag följer kärleken . Åh ... Jag är inte ... 
Smickra inte dig själv . 
Nu när vi hjälper till , kanske ni har en chans . 
Du vet . En liten chans åtminstone . 
Vi rensar ytterdörren . 
- Hallå ! - Vill ni tävla ? 
Okej , det är lugnt . 
Scanlans hand Är du säker på det här ? 
Jag har aldrig gjort en plan förut . 
Ingen annan i gruppen heller . 
Vi är körda hursomhelst . 
De är inne . 
Tillbaka till de andra . 
Se upp ! 
Keyleth , få ner mig dit ! 
Nej , nej ! 
Raishan ? 
Vad gör hon ... 
Spring ! Det är instabilt ! 
Håll er nära ! 
Jag såg Raishan och hon hjälpte inte till . 
Hon slåss åtminstone inte mot oss . 
Jag ogillar det . 
Inkommande ! 
Här borta , fulis ! 
Vad blir det till middag ? 
Jag önskar att du kunde ta saker lite mer på allvar . 
Det är inte bra . 
Täcker du mig ? 
Ja . Var försiktig . 
Bära eller brista . 
Åh , det sved ! 
Kom igen , bjässen ! 
Det räcker ! 
Kash ! 
Vänta . 
Är det ... Nej ! 
Herregud , nej ! 
Titta inte . 
Kash ! 
Vax , vi drar . 
Kom ! 
Shaun . Få bort Zahra härifrån . 
Du då ? 
Han har förstört för många liv . 
Vi avslutar det här . 
Lycka till , din snygga dåre . 
Kash , jag förstår inte ... Han ska inte dö förgäves ! 
Raishan sa väl att själsankaret är Thordaks kraftkälla ? 
Så hur träffar vi det ? 
Kiki , redo för den stora ? 
Ja , för fan ! 
Nu ! 
Är du okej ? 
Fungerade det ? 
Det är omöjligt . 
Det måste ha hänt något . 
Vi stannar inte för att ta reda på det . 
Kom igen , snälla ! 
Fan ! Jag trodde att jag hade det ! 
Bäst att du löser det . 
Zahra , jag kan inte . 
Till och med när jag tvekade , så visste Kash att reliken var menad för dig . 
Thordak har tagit så mycket . 
Låt den jäveln blöda för det . 
Scan-man ! Jag har hittat ett ! 
Du får nog räkna om , kompis . 
Okej . Bäst att vi förstör dem fort innan de tar över . 
Vänta , det känns fel . 
De är väl bebisar ? 
Driver du med mig ? 
Vi kanske ska vänta tills de är lite äldre ... 
Grog , det är dåliga ägg . Hör du mig ? 
Gör omelett till mig , för helvete ! 
Var det ... Var det för mycket ? 
Raseri ! 
Lite rädd , lite upphetsad . 
Nej ! Överallt utom ansiktet . 
Kukblixt ! 
Åh , nej . Gör inte så . 
Vart fan ska han ? 
Grog och Scanlan måste väl ha lämnat nästet ? 
Det är inte så vår tur fungerar . 
Kom igen ! Fy tyst på dem ! 
Nej , stopp , stopp . 
Det är jag ! 
Oj , du ser för jävlig ut , kompis . 
Jag känner mig så också . 
Vi måste sticka innan ... 
Jävlar , göm dig ! 
Mitt blod ! 
Mina arvingar ! 
Nej ! 
Du , du har varit plankillen idag . 
Har du en till ? Va , jag ? 
Jag slår bara på saker . 
Vänta . 
Jag slår på saker . 
Vem gjorde det här ? 
Ja . Det var jag . Jag gjorde det . 
Förlåt , jag trodde att det var äggbuffé . 
Mina barn föds så hungriga . 
Ditt svedda kött kommer att fylla deras magar som kompensation . 
Jaså ? Hur ska de äta mig med ett tak på sina huvuden ? 
Dåre , du vet inte vad du gör ! 
Det gör jag aldrig . 
Du trotsar en kung ! 
Helvete ! 
Vi dör . Vi dör nu ! 
Utgången . 
Scanlan ! 
Jösses ! Vilken åktur ! 
Eller hur , Scanlan ? 
Scanlan ? 
Vakna . 
Nej . 
Kan ... Kan du fixa honom ? 
Fan ! 
Snälla ... Du måste fixa honom . 
Mina barn . 
Vårt herravälde . 
Min värdefulla framtid . 
Förstörd ! 
Jag ska avlägsna ert kött ! 
Vax , vad gör vi ? 
Vi gör en sista insats . 
Pike ! Vänta ! 
Lita inte på någon annan än dig själv . 
Det är inte rustningen . 
Det är jag ! 
Jag är här , Thordak . 
Din jävla förrädare . 
Raishan . 
Utplåna vår fiende . 
På din befallning , min kung . 
Din bitch ! 
Hur vågar du ? 
Jag frigav dig . Följde dig . 
Satte ihop din konklav . 
Du skulle ha hållit ditt ord . 
Smaka på min sjukdom . 
Nåväl . 
Jag återkommer . 
Vex , Vax . 
Den här världen kan vara ond . 
Fylld av de som vill förstöra den . 
Men den flödar även av hopp . 
Ta hand om varandra , skydda era vänner ... Och kom ihåg ... Inget är starkare än kärlek . 
Thordak ! 
Nej . 
Jag vill ha ont ett tag . 
Han är vid liv men ... Han vaknar inte . 
Men han kommer väl ... - Eller hur ? - Jag vet inte . 
- Vi gjorde vårt bästa . 
- Men det får inte tillbaka dem . 
Mor . Percy . 
Gå till henne , bror . 
Jag hade fel om Raishan . 
Det kvittar . 
Det gör det inte . 
Förlåt , Vax . 
Jag ska säga det till henne med . 
Vad gör du ? 
Beundrar vad vi lyckades åstadkomma , tillsammans . 
Jag ... Jag vill tacka dig för att du hjälpte oss i konklaven . 
Ditt tack behövs inte . 
Vi hade båda anledning att hata Thordak . 
Din allians var ändå uppskattad . 
Vad händer nu för Vox Machina ? 
Svårt att säga . 
Jag vet inte hur vi ska kunna fortsätta som vanligt . 
Vad ska du göra ? 
Vad jag än önskar . 
Är det ... Vänta , vad är det ? 
Din instinkt är korrekt , tjejen . 
Jag har alltid tyckt att du är den smarta , Keyleth . 
Släpp aldrig garden runt din fiende . 
Du gav mig exakt vad jag behövde . 
Rör dig inte ! 
Kom ni för att gratulera mig ? 
Vi har redan dödat en drake idag . 
Vi kan döda två . 
Vilket övermod ! 
Men jag ska säga tack . 
Jag hade inte kunnat göra detta utan Vox Machina . 
Och inte det som kommer . 
Fan ! 
Vart tog hon honom ? 
Är du okej ? 
Inget är okej . 
