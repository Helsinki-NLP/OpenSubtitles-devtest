Alice . 
Även om jag inte är här finns jag alltid med dig . 
Oavsett vad som händer , vakar jag alltid över dig . 
Houston . Det här är Birdsong . 
De lever . 
Jag måste ha svimmat av . De andas . 
Jag kan se deras andedräkt ! 
Men de var döda ... Herregud ! 
Jag kan se deras andetag . 
De lever . 
... svimmat av . 
De andas . 
Jag kan se deras andetag . 
De lever . 
De andas . Jag kan se deras andetag . 
Sätt dig , pappa . 
Sätt dig . 
Hör på . Mamma är död . 
Jag är ledsen . 
Hon dog i olyckan . Ursäkta ? 
Hennes kropp är kvar där uppe . 
Du tillbringade just två dagar med henne i stugan . 
Jag hörde det . 
Mamma lever . Hon är bara inte med oss . 
Vi miste vår mamma . 
Och det finns en annan Alice . 
Det är hennes mamma som kom tillbaka . 
Det finns nån annanstans . 
Det har nåt med CAL att göra . 
Mamma har en mentalsjukdom . 
Vad hon än har sagt , är det inte sant . 
Mamma lever . 
Du har fel , pappa . 
Det är nåt fel på maskinen . Bilden är förvanskad . 
Visa mig . 
Anklagelserna är att mr Caldera sköt befälhavare Paul Lancaster på 60556 Lexington Avenue cirka kl 21 : 05 måndagen 8 november 2021 . Dessutom att mr Caldera kastade mr Ian Rogers från aktern på SS Bernice , utanför Santa Barbaras kust kl 23 : 35 söndagen 17 oktober 2021 , vilket orsakade att mr Rogers drunknade . 
Fortsätt . 
Mr Caldera säger att han inte är personen som begick dessa brott . 
Dessutom begär han ett polygraftest för att bekräfta hans identitet och minnet av dessa saker . 
Ni måste jämföra mitt DNA med invånaren av Bud Calderas lägenhet . 
Men ni förnekar inte att ni är Henry Caldera . 
Vi har nog redan fastställt att den jag inte är , är Bud Caldera , så kallad . 
Vad jag skulle påstå är att dessa två herrar är samma person . 
Med all respekt , det är de inte . 
Ni måste fastställa var Bud Caldera bor och vad hans personliga och ekonomiska omständigheter är . 
Kortfattat , jag behöver hjälp att ta reda på vad hans liv är . 
Läs den här . 
Gud vet vad den kostade . Förmodligen miljoner . 
Men hon har tagit en satans yxa och gett den 40 jävla hugg . 
Jag beklagar . 
Å Europeiska rymdbyråns vägnar . 
Hon får behandling . Vi kommer att avskeda henne . 
- Jaså ? - Ja . 
Jag minns 1964 , den första intagningen av kvinnliga astronauter . 
De hade just genomgått sin fysundersökning , och Steven Winderuss , verksamhetschef på den tiden , skrev en rapport angående problemet med kvinnor i rymden och krångligheterna med att matcha ett temperamentsfullt psykofysiologiskt objekt t.ex. en kvinna , med en komplicerad maskin , t.ex. en rymdfarkost . 
Det är ... ett problem vi aldrig löst . 
Henry , är du inte bekymrad över det här ? Nej . Nej . Vadå ? Det är ett föremål . Vi har liv att leva . 
Vad ... Vad är det som händer ? 
Varför är jag inlåst ? 
Varför är jag här ? 
Talar du engelska ? Talar du ryska ? Vänta , vänta , vänta ! Snälla ! Vänta . Vänta , snälla ! Hallå ? Snälla , kom tillbaka ! Snälla ! 
Har hon sin telefon ? Jag vet inte . 
Varför vet du inte ? 
Jag måste prata med henne om några saker . 
Du trodde ju att hon var död . 
Alice . Ät din frukost . 
- Den smakar som skit . 
- Den smakar inte som skit . Du har aldrig smakat skit . 
Du får inte träffa din mamma om du tror på allt skräp hon säger . 
Det här är inte PTSD . Det är inte psykos . Det är inte schizofreni . 
Det är vad alla med schizofreni och psykos säger . 
Jag måste hem till min dotter . 
Du spelar väl piano ? 
Spela . 
Det bröt ut en brand i min stuga . 
Innan dess såg jag min dotter . Den riktiga . Jag har inte sett henne sen innan jag åkte till rymden . 
Spela . 
Är du mamma ? 
Du reste med din dotter . 
Hon var väldigt sjuk efter branden , men nu mår hon bra . 
Hon är med sin far . 
Jag kunde lukta henne . 
Den riktiga Alice . 
Jag ... Jag kunde känna doften av min dotter . Jag ... Om det här tillståndet inte behandlas kommer det att bli värre , tro mig . 
Varför förhindrar ni mig från att träffa henne ? 
Snälla . Hon är min älskling . 
Hon är min älskling och jag har förlorat henne . 
Du är gravid . 
Du vet att vi måste ta ett graviditetsprov innan vi ger litium . 
Det kan vara giftigt för fostret . Vad ? 
- Normalt skulle vi ge dig ... - Åh , nej . ... 1 800 milligram litium-7 för att dämpa dina symptom , men du är gravid i ett tidigt skede . Fjärde veckan . 
Vi har utformat en alternativ läkemedelsbehandling åt dig , men du måste åta dig att genomföra den . Annars måste vi chocka dig igen . 
Jag kan inte föda barnet . 
Om jag föder barnet , hur ska jag ta mig tillbaka till henne ? 
Snälla . Ta de här tabletterna . 
Jag ser att du har ont . 
Jag kan hantera smärta ! 
Det här är inte vansinne . 
Jag måste återvända till henne . Förstår du ? Jag kan inte vara här . 
Vad fan är det för oväsen ? 
Det finns en annan gäst . 
Du kommer inte att se dem . 
Obotlig . 
Snälla , gå inte ... 
Det är ... Det är du . 
Det är flammor ... Eld ! Eld ! 
Kapseln brinner . Fyrtio . Fyrtiotvå . 
Det är hett . 
Hett . Världen är uppochnervänd . 
Det är Irena . Jag måste träffa dig . Det är brådskande . 
Har ni nånsin träffat Ian Rogers ? 
Jag vet inte vem det är . 
Har ni nånsin varit ombord på SS Bernice ? 
Inte vad jag vet . 
Träffade ni Paul Lancaster ? i ert hem i East Hollywood ? 
Jag har inget hem i East Hollywood , därför träffade jag inte Paul Lancaster . 
Har ni nånsin träffat Paul Lancaster ? 
Många gånger . 
Under vilka omständigheter ? 
Jag minns inte de ursprungliga omständigheterna , men vi var båda anställda av NASA och arbetade med ISS-programmet : jag som chefstekniker på Raketdriftslaboratoriet , han som astronaut och missionsbefälhavare . 
Sköt ni Paul Lancaster ? Nej . 
Men jag kan nog ha dödat honom . Hur ? 
Jag uppfann en maskin som orsakade eller snarare möjliggjorde , en dödlig olycka i rymden . 
När trollmor har lagt ... Jag vill gärna höra dig spela . 
- Hej ! 
Bad ... Bad de dig komma ? 
Har du ... Har du pratat med Magnus ? 
Träffade du Alice ? 
Jag har ställt många frågor om den här åkomman . 
Varför spelar du inte ? 
Jag har aldrig hört dig spela piano förut . 
Ilja , det här kan låta galet , men det ... det är ingen åkomma . 
Hör på , jag har läst om Henrys arbete . 
Vet du var Henry Caldera är ? 
Vad han gör ? Kanske jag kan prata med honom . 
De kallar det " astronaututbränning " . 
En känsla av dissociation . Paranoia . En känsla av att bekanta platser och människor är bedragare . 
Det har hänt många gånger . 
Den goda nyheten är att de kan medicinera det . 
Varför har du kommit hit ? 
Irena är sjuk . Hon hoppas att jag ska ta över . 
Det måste finnas nån här som kan ta hand om folk . 
Ilja , jag har hört inspelningar av radiosändningarna från hennes kapsel . Den upplöstes i rymden . Hon dog . 
Irena var kroppen som kolliderade med ISS . 
Paul dog inte . Det var jag . 
Jo , om hon kolliderade med ISS , hur kan hon vara här ? 
På samma sätt som jag är här . 
Vi k ... Vi kom ... från nån annanstans . 
Den enklaste förklaringen på att ni båda är här är att ni båda återvände levande . 
Jag minns inte henne . 
Hon är chef för Roskosmos , och jag minns inte henne . 
Jag minns inte CAL . Jag minns inte Henry Caldera . Jag minns inte min dotter . 
Så det är nåt fel med ditt minne . 
Försvinn . 
Det finns så mycket för dig här , Jo . 
Sluta sörja och bli bättre . 
Snälla . 
Om du inte blir bättre , blir du bara sämre . 
Jag trodde jag såg henne . I snön . 
Och för ett ögonblick blev jag ... Jag blev så glad att se henne igen . 
Jag kände hur mycket jag saknade henne och hur mycket jag älskade henne och hur ledsen jag var . 
Och sen var hon borta . 
Jag är fast i mitten . Och de går båda igenom saker som jag inte har nån aning om . 
De har hemligheter som jag inte är en del av . 
Jag vet inte hur jag ska gå vidare från det . 
Eller hur jag ska få Alice att gå vidare från det . 
Hur ... Hur kan vi återförenas igen ? 
Vill du återförenas igen ? 
Det känns som om vi alla svävar i rymden . 
Det känns bara som om vi alla svävar i rymden . 
Jisses , det må jag säga , - det här är bättre än jag är van vid . - Henry . 
Du får mig att känna mig märkligt bättre . 
Vad ? 
Vad är annorlunda ? Kom . 
Du vet , för länge sen , när jag genomgick utbildning , åkte Irena Lysenko upp i rymden . Och ... Och hon kom ner igen välbehållen . 
Och jisses . Åh , vilken snygg tjej hon var . 
Jag träffade henne aldrig . Men sen åkte jag iväg . 
En lång tid var jag inte mig själv . 
Men det är då jag minns att jag hörde att det skedde en olycka där uppe och att Irena Valentina Lysenko faktiskt kvävdes till döds . 
Det är sjukdomen som får dig att tro det . 
Henry , vi genomgick båda en olycka . Det kändes märkligt att komma tillbaka . Det var det fanimej . 
Du sa att du kände en annan person gå vid sidan om dig . 
Nån har sovit i min säng och burit mina kläder och ätit min satans gröt . 
Du är experten . Om jag börjar ta de här igen , kommer det att jämna ut min lilla personlighetsstörning ? 
Henry , vad är det med dig ? 
Jag är inte Henry . 
Henry är borta . 
Och peppar , peppar , om jag har tur , så kommer han aldrig tillbaka . Men han kommer att minnas vem han var , och han kommer att leva min ålderdom , mina beroenden och mina jävla misslyckanden . 
Du måste följa med mig till St . Sergius . Jag kan hjälpa dig . Jag behöver inte hjälp . 
Jag ... Jag är killen som vann Nobelpriset . 
Jag blev fotograferad med Reagan och Muhammad jävla Ali . 
Det är jag . 
Och du kan fortsätta att förneka och mörka det som du alltid har gjort . 
Tror du på spöken ? 
Jag vet inte . 
Ibland tror jag att min pappa är här . 
Jag vet att han dog , men ibland tror jag att han är här . 
Wendy , jag ... jag tror att min mamma är död och att det finns en annan som lever . 
Jag skulle byta plats med dig . 
Hälften levande och hälften död är bättre än helt död . 
Kanske en del människor kan finnas där och inte finnas där . 
Vad hände med din pappa ? 
Han var lite galen på mammas begravning . 
Jag vet inte . 
Han åkte för att träffa en astronaut och blev skjuten . 
Han är på sjukhuset nu . 
Jag är lite ledsen . 
Jag är fortfarande ledsen över min mamma . 
Jag tror att jag såg hennes spöke . 
Men din pappa är cool . 
Han är tjurig . 
Han är en snäll pappa . 
Ja . Jag antar det . 
Pappa , jag vet att det är påhittat det hon sa . 
Jag vet att hon inte dog . 
Det gläder mig att höra . 
Så , kan vi åka och träffa henne ? 
- Vill du ha grejorna i lådan ? 
Några saker de hittade utanför stugan Ja . 
Alice , sista chansen . Vill du kolla att du inte har lämnat nåt där uppe ? 
Kan du höra mig ? 
Vill du leka en lek ? 
Är mamma där ? 
Jag vill veta om jag verkligen såg henne vid stugan . 
Snälla ? 
Jag vill prata med henne . Snälla . 
Vi ska åka nu . 
Så där . 
Jag ska sluta leta efter mamma . 
Det finns en annan Alice . Hon finns på ett annat ställe . 
Hon fick mamma i stället för mig . 
Det är en bra inställning . 
Jag kan inte vara arg på andra Alice bara för att hon hade mer tur . 
Jag är väldigt stolt över dig . 
Är jag modig ? 
Du är otroligt modig . 
Och polygrafen ? 
Du klarade det med glans . 
Och DNA-provet ? 
Om jag har rätt , så vrider sig mitt i en annan riktning än det ni hittade hemma hos Bud Caldera . 
Nix . DNA:t är exakt detsamma . 
Och polygrafen bevisar bara att du tror att det du säger är sant . 
Det är sant . 
Sanningen är en bristvara nuförtiden . 
Har det gått er förbi ? 
BERNICON IV . GÄSTLISTA Henry , även känd som Bud Caldera , Jag anklagar dig formellt för mordet på Ian Rogers och mordförsöket på befälhavare Paul Lancaster . 
Ni har rätt att tiga , men det kan skada ert försvar om ni inte nämner under förhör något ni senare förlitar er på under rättegång . 
Då går vi vidare till kvällen för den så kallade " dubbla händelsen " . Tre veckor efter mordet på Annie Chapman , 30 september 1888 . 
Det var en blöt , eländig kväll . Och oerhört mörkt . 
Kl 01 : 00 styrde klubbens förvaltare sin häst och kärra genom valvet där in i passagen . 
Hästen hoppade åt vänster , skrämd av nåt som lurade i grändens skuggor . 
Jack Uppskäraren . 
Om vi går vidare till nästa plats , kan jag visa er var . 
Vad i helvete ? 
Jag är pensionerad polis . 
Jag vet . 
Lev ditt bästa liv , Ian Rogers . 
Hur mår du ? 
Vilka är männen där uppe ? Det finns bara en man . 
Vem är han ? 
Den första mannen i rymden . 
- Vad ? 
- Ta din medicin . 
Spela på pianot . 
Gör saker din kropp är van vid . Det hjälper . 
Annars kommer du att brista , tro mig . 
Dog jag där uppe ? 
Kan jag ta mig tillbaka ? 
Kan jag nånsin ta mig tillbaka ? 
Finns det två av dig ? 
En död , en levande ? 
Finns det två av mig ? 
Hur förbättrar det vår vetskap om oss själva ? 
Men om det här är vad som händer där uppe ... Nu räcker det . 
Du har ett barn här att vara mamma till . 
Och kanske ännu ett på väg . 
Acceptera det här och släpp taget . 
Hur skulle jag kunna det ? Jag ... jag ... jag kan inte . 
För vad det än är , så kan det inte göras ogjort . 
Du kan inte ändra på det . 
Nånsin . 
Det är gjort . 
Lev . 
Jag har tänkt på den andra Alice . 
Jag tror att hon känner att det är okej . Att du är här med mig . 
Jag känner att hon tycker att det är okej . 
Vi förlorade båda nån , men vi fann båda nån också . 
Det betyder inte att vi måste glömma den andra . 
Bara att vi måste acceptera det . 
Accepterar vi det ? 
Du är en enastående ung människa , Alice . 
Din mamma skulle vara otroligt stolt över dig . 
Är du stolt över mig ? 
Jag behöver en mamma . 
Jag behöver en Alice . 
Det är jag . Mamma , det kan vara jag . 
Det här är vad jag såg . 
Det här är vad som kolliderade med ISS . 
Alice ritade det här . 
VALJAN Hon hörde förmodligen dig prata om det . 
Jag försöker vara rationell , Magnus . Min man är här . 
Min dotter är här . 
Det är uppenbarligen samma värld som jag lämnade . 
Men vad ? 
Jag ska börja ta tabletterna om det betyder att jag ... Att jag slipper leva på den här knivseggen . 
Och det här barnet ? 
Du ville ju alltid ha ett till , men vi har inte pratat om det sen din rymdfärd . 
Är vi i skick att ta emot det ? 
Vill du ha det ? 
Vill du ? 
Mitt namn är Irena Valentina Lysenko . 
Jag är verkställande chef på Roskosmos . 
TILL : UTSKICKSLISTA ASTRONAUTER År 1967 blev jag den andra kvinnan i rymden . 
Sen den gången under Sovjetunionen , och sen kommunismens fall , har det varit min börda och mitt ansvar att dölja ett enkelt faktum om rymdresande . 
Att det driver folk till vansinne . 
Vi vet det här . 
Ni vet det här . 
Vi låtsas att det inte är sant , men väldigt många av oss ser och hör saker som inte kan förklaras kanske inte ens genom att kalla det " vansinne " . 
Jag undrar om ni kanske vore villiga att rapportera några av era egna problem anonymt till mig . 
Paul , släpp . 
- Jag ser nåt ! 
Jag är ledsen . 
Saker är annorlunda . 
Magnus , verkar ... verkar jag som din Jo ? 
Jag älskar dig . 
Jag älskar dig och jag ... Jag vill ha dig mer än jag ville . 
Jag också . 
Får jag sitta hos dig ? Visst . 
Tack för att du tog hand om henne . 
Här . 
- Vad heter du ? 
- Irena Valentina Lysenko . 
Men mina vänner kallar mig Valja . 
Ner i kaninhålet med dig , Alice . 
Mot oändligheten och vidare ! 
Ge mig bara en minut , okej ? 
Mamma ? 
Får jag fråga dig en sak ? 
Om det som hände hände om jag är härifrån och pappa är härifrån och du är därifrån var kommer babyn att vara ifrån ? 
Alice , även om jag inte är här så finns jag alltid hos dig och pappa . 
Du förstår nog inte hur mycket jag ... Jag ville bara finnas där och se dig växa upp . 
Oavsett vad som händer kommer jag alltid att vaka över dig . 
Och mitt hjärta slår med dig , älskling . 
Jag älskar dig så mycket . Mer än du nånsin kan föreställa dig . 
Min älskling . 
