TIDIGARE I SERIEN ... 
Du får göra om den . 
Stirling , karlen som du grillade på gårdagens fest . 
Den där bysten du gjorde , kan du lära mig göra en ny ? 
- Ge den tillbaka ! - Vill du ha den ? 
- Kom och ta den ! - Ge mig min bräda ! 
- Du kan inte ens köra . 
- Du ska få se . 
- Bort från min bil ! - Kör ! 
Du skulle bara våga ! 
Ta det lugnt . 
Du kör för fort . 
- Sväng ! - Jag försöker ! 
- Försök hårdare ! 
Jag vill ha en ny bil . 
- Varför ? 
- För att hålla henne borta . Mia . 
Någon måste ta kontroll över familjen , så nu flyttar jag in . 
Jag vill träffa Mia . 
Hon behöver mig . 
Någon dog på grund av elavbrottet . 
Wayne vill att jag håller det ifrån tidningarna . 
Jag vill att vi arbetar ihop . 
Får jag fem minuter med honom , får jag honom att investera . 
Murray Doull . 
- Gäller ditt erbjudande ännu ? 
- Ja . 
Kvinnor åker inte till rymden längre . 
Bättre att bli skönhetsdrottning , va ? 
Åttio Mississippi , 79 Mississippi , 78 Mississippi , 77 Mississippi , 76 Mississippi , 75 Mississippi , 74 Mississippi . 
Jag mår bra . 
Du verkar inte må bra . 
- Krocken , Tilly ! Det ... 
- Det är över . Du är okej ... 
Det är inte okej . Vi måste betala de där arslena för deras usla bil . 
Tusen dollar . 
Och de ville göra mig illa . 
De kom efter mig på min strand . 
- Det är fortfarande din strand . 
- Nej , stranden är deras . 
Trettiotre Mississippi , 32 Mississippi , - 31 ... Skylab ! - Trettioett ... 
Skylab ! 
Åh , det är tidigt . 
Syns den bättre ? 
Den är närmare . 
Tänk om någon ser vagnen gunga och tittar in ? 
Det är det 17:e tillägget i australiska konstitutionen . " Om vagnen vajar , kom inte och knacka . " 
Konstitutionen . Den har aldrig gjort något för mig . 
Är jag " bra Sandy " eller " dålig Sandy " ? 
- Min farsa är en idiot . 
- Det är klart . Han är polis . 
Du känner inte till hälften . 
Vänta ! Är det Rocco ? 
Var inte rädd , han kommer inte hit . 
Han kunde inte bry sig mindre . 
Ja . 
Killar som jag har mördats för mindre . 
Vi ses . 
Du är en väldigt , väldigt " bra Sandy " . 
Vad är klockan ? 
Sju . 
Hela gatan vaknar upp . 
Är du vaken ? 
Du var ute . 
Jag behövde träffa Jude . 
Varför ? 
Kvinnosaker . 
Lämna mig ifred . 
ELSTREJKER KAN DRABBA INFRASTRUKTREN 
Francesca , du är en romersk gudinna . 
Alltså ... 
Francesca tror inte att Kanal Sju:s nyheter vet om dödsfallet på sjukhuset . 
- Tror inte ? 
- Vi får veta ikväll klockan sex . 
Om de vet om det , och du inte ... och Wayne inte står till svars ... 
I så fall blir vi slaktade . 
Jag har inte sett dig i slips på länge . 
Man behöver ingen på barrikaderna . 
Det är synd . 
Den klär dig . 
I slips kunde du ha fått en bättre deal . 
- Du erbjöd mig ingen deal . - Ja , okej . 
Jag har ingen aning om vad ni vill . 
Gazza och hans kompisar bara förhalar . 
Hur skulle det vara med garantier för ett år , och tio procents lönesänkning ? 
Är det garantierna eller lönen ? 
Gazza säger att det är båda . Men det är alltid pengarna i fickan . 
Är det ? 
Hur skulle det vara med jobb garanterade för ett år , och fem procents lönesänkning , exklusive , 
nej , inklusive övertid ? 
Vi har en deal . 
Dag ett med Bissett Star Broadcasting ! 
Jag kanske hade haft det bättre på den döende strömförsörjningsfirman . 
Det är bara en enkel omfördelning av tillgångarna . 
Mercan mot skåpbil och utrustning . 
Låter inte kanon . 
Vi har Barrys nya skåpbil , verksamheten växer fort . 
Så som du ofta gillar att påpeka , inga barn , ingen fru . 
Vad skulle jag annars riskera ? 
Varför måste jag ha snaran om halsen ? 
Miss Universum ? 
En intervju med grundaren av " den döende strömförsörjningsfirman " . 
- Nej . 
- Jo . 
Mia ! 
Skola . 
Mia ! 
- Ord ? 
- Jag går ingenstans . 
Jag träffar ingen . Skolan . Stranden . Inget . 
Kom igen . 
Det har gått flera dagar . 
Mia ! 
Kan du en gång lämna mig i fred och oroa dig för Tilly . 
Hon är besatt av Skylab och har gett upp hoppet om att vara första kvinnan på Jupiter ! 
- Tilly ? 
Vad ? - Har du inte märkt ? 
Okej , jag ska prata med henne . 
Skola . 
Jag skojar inte , Mia ! 
Stig upp ! 
Jösses . 
James Stirling ? 
På allvar ? 
Det är Yellagonga . 
Era män kallade honom kung , men han var ledaren av Wahdjuk Noongar under kolonins första tid . 
Bilya . 
Han är en legend för vårt folk . 
Han förtjänar att bli hyllad , inte Stirling . 
Jag ber om ursäkt , mr Williamson . 
Bilya , du är här för att lyssna och lära dig . Inte föreläsa . 
Imponerande entusiasm , Bilya , men jag tror din lektion börjar . 
Jag ber om ursäkt . 
Han lär sig . 
Han är ung . 
Men du ... du tycks ha en god förståelse för vår historia , Eileen . 
Du borde vara på radion . 
Vi har erbjudits några intervjuer för lokala lärare , att prata om vår historia och deras arbete . 
Det kommer att höras långt , kanske i hela delstaten . 
Jag vet inte . 
Det är en chans för en lärare från ursprungsbefolkningen att visa vilka framsteg vi gjort under de gånga 150 åren . 
Okej . 
Låter bra . 
- Jag måste gå på lektion . 
- Okej . Tack , Eileen . 
Skit , Francesca , vad är det nu ? 
Har du gjort av med fler , va ? 
Vi har en plan . 
En deal att få slut på strejken och hålla företaget i gång . 
Att få företaget att växa . 
Vi har förstått att fackföreningarna godkänner en fem procents lönesänkning . 
Tillsammans med inbesparingar som vi gör med leverantörer och processer , betyder det att vi kan få slut på strejken - och gå vidare . 
- Men jag måste acceptera det . 
Vi rekommenderar att du gör det . 
Det är en bra deal , Wayne . 
Ni tror väl inte att jag läser allt detta , va ? 
Jäklar ! 
Hur ser jag ut , Frannie ? 
Jag tänker planka in på farsans tv-intervju och vill se bra ut . 
Du är jättesnygg . 
Om du inte har tid att läsa , kan vi sammanfatta det åt dig . 
Jag vet ändå att det är skit . 
Jag hoppas du tar det lugnt med mig , det är inte mitt företag längre . 
- Nej , inte officiellt . 
- Oroa dig inte , mr Doull . 
- Jag ska vara snäll . 
- Får vi göra er sällskap ? 
Wayne . Vilken trevlig överraskning . 
Kul att se dig , Tony . 
Du kan inte hållas borta , va , pappa ? 
Och du , min son , kan inte motstå en kamera . 
Jag tänkte ni kunde ha användning för ett vackert ansikte . 
Familjen Doull har alltid varit ledare , särskilt under tuffa tider för Perth . Wayne fortsätter den traditionen . 
Och hur stolt är du över din sons insatser under dessa svåra månader , sedan han tagit över ? 
Mycket stolt . 
Jag är säker på att det finns en lösning . 
Tack vare Waynes hårda arbete och hans nya vackra chef Jude . 
- Du är inte David Frost precis . - Håll käft . 
Ska jag prata ? Okej . 
Jag har pratat med fackföreningen och är ganska säker på att jag förstår deras behov och önskemål . 
Vi fokuserar förstås på hur företaget ska gå framåt . 
För att vara hållbara fokuserar vi på långsiktig sysselsättning . 
Jag tror att vi hittar en kompromiss som löser det . 
Där har vi ett smutsigt ord ! " Kompromiss " . 
Dessa giriga fackföreningar måste förstå att detta företag , detta anspråkslösa familjeföretag ... 
Ett familjeföretag som behandlar sina anställda som familj . 
Alltid gjort det , kommer alltid att göra . 
Ja , jag kan gå i god för Murray . 
Jag har jobbat på detta företag i nästan två årtionden . 
Jag han känt Murray nästan lika länge som min man . 
Platsen känns faktiskt som familj . 
Tills du avskedade din man . 
Kanske vi klipper bort det ? 
Inget illa menat , Tone . 
Du blev uppsagd , du fick inte sparken . 
Det är okej , Wayne . 
Men du kan väl berätta för kameran , hur det känns för din lilla , lyckliga strömfamilj att ha orsakat sorg i en annan familj ? 
Vad pratar du om ? 
Mr Doull , under din sons ledarskap , har dispyten lett till ett dödsfall på Scarborough Beach Sjukhus . Det rådde brist på företagets delar som de hade behövt för att få igång sin nödgenerator . 
- Vad ? 
Ett dödsfall ? 
- Vi måste sluta nu . 
- Ja . - Har du blod på händerna , Wayne ? 
- Hej ! - Mick , det räcker . 
Fan ta det här . 
Kassett - och batteribyte . 
Ursäkta . 
Tony . 
- Kan du hjälpa honom ? 
- Ja . 
Ni sänder inte det där . 
Den tappre är taktfull , mr Doull . 
Tappre ? 
Plötsligt anklagad för korporativt dråp . 
Men det är väl det som du kallar " story " ? 
Något i den stilen . 
Och något i den stilen är välbetalt ? 
Det är tanken . 
Jaha ... 
Jag börjar förstå mig på din verksamhet . 
Vi borde äta lunch ihop ... tillsammans med våra damer och diskutera allt detta . 
Utmärkt idé , Murray . 
VAR GOD RING 
Det är avgångsvederlag . 
Alltså ... 
- Det var en överraskning . 
- Jag försöker bygga något . 
Allt du gjorde idag var skada . 
Jag trodde att vi skulle ta upp Miss Universum , - inte jävlarna som gav mig sparken ! 
- Du , vi tar upp all möjlig skit som vi kanske inte gillar . 
Kan du inte hålla tyst i en timme eller två ? Är det omöjligt ? 
Jag är ledsen , Mick . 
Verkligen . 
Ja ... Du är min bror , och därför kommer det inte att funka . 
En till dag som denna och jag förlorar mitt jobb . 
- Mick ... 
- Jag också . 
Inget illa menat . 
Snälla . 
Behåll dem . 
Nej , fan . 
Jag måste betala för en krockad bil . 
Fan ! 
Nu räcker det . 
Kom igen . 
- Varsågod . 
- Tack . 
Vilka vågor ! 
Efter London kändes de som liv . 
Även under de mörkaste perioderna , kunde jag gå dit . 
Och fly världen , bara för några sekunder . 
Vågorna var dina , du kunde göra vad som helst . 
Det kan du fortfarande . 
Stranden ... De där killarna är där . 
Mia , åt fanders med dem ! 
Nu kan vi antingen vända om , och vara tillbaka vid tedags , eller så kan vi få din bräda fixad . 
Varför kallas han " Spindeln " ? 
Han klamrar sig fast vid brädan , man kan inte skaka loss honom . 
Han faller aldrig . Han är lite som du . 
Ser man på ! 
- Bobby Foden ! 
- Goddag , Gerald . 
Fem fan är " Gerald " ? 
Det är det största hedersmärket som jag någonsin sett . 
Den som gör så mot en bräda är ett arsle . 
Om de inte gillar dig , betyder det att du är ett anti-arsle . 
Vilket betyder att du är min typ . 
Jag vet att du kan fixa den . 
Jag vet inte om jag borde . Jag menar det . 
Det är en del av brädans historia . 
- Det är en del ... - Mia . ... av Mias historia . 
Fint namn , Mia . 
Jag vill bara få bort det så fort som möjligt . 
Du gillar stora vintervågor , va ? 
Det är väl klart ? 
Säg mig har snubben fortfarande min husvagn ? 
- Din husvagn ? 
- Ja . Han vann den i skumt kortspel . 
- Vill du spela för vagnen igen ? 
- Nej . 
Titta var jag hamnade , du din jävel . 
Kom . Nu tar vi bort vaxet . 
Tack , mrs Doull . 
Det var härligt . 
Tack för att ni visade mig hur stiligt livet är här . 
Det är klart att Mick också har visat mig . 
Hans videoklipp om staden och tävlingen är så filmiska ! 
På tal om det , har ni båda biljetter - till miss Universum-finalen ? 
- Ja , naturligtvis . 
Då ska vi få er backstage innan det börjar ! 
Om ni vill , så klart . 
Du vet hur man väljer dem , Mick . 
Det gör jag också . 
Jag gillar din verksamhet . 
Det kommer att finnas mer av allt på 80-talet . 
Mer tv , fler kanaler , fler kändisar . 
Det är vad folk vill ha . 
Jag ger dig 150 000 , för 49 procent av firman . 
Det är inte en 300 000 dollar business , Murray . 
Det vet du . 
Du vet också vad det här kan bli . 
Och vad det kan erbjuda på vägen . 
Titta på den här fantastiska hamnen . 
Om jag bodde i Australien skulle jag vara här varje dag . 
Jag ger dig 150 000 , för 40 procent av firman . 
Trettio procent . 
Och kassetten från idag . 
Okej . 
Trodde jag skulle säga sanningen . Ja . 
Men inte om du då blir avstängd eller jag sparkad . 
- Morbror Adam varnade mig . 
- Vad ? 
Vad varnade han om ? 
- Att du bockar för dem . 
- För att behålla mitt jobb . 
För att behålla vårt hem . 
Det är lätt för honom ... 
Gå in . 
MARK , INTE ALLMOSOR ! Ni tror att klistermärken ändrar världen . 
STULEN MARK BEFRIA SVARTA AUSTRALIEN 
Fem , fyra , tre , två , ett och stopp . 
Hur gick det ? 
Kom igen , Till . Du bad om testet . 
Du måste vara självsäker . 
Jag vet inte , sekreterarskolor vill ha 100 ord per minut ... 
Ja , men jag tror att de vill ha dem i rätt ordning . 
Jag beundrar att du har mer realistiska mål än att åka till månen . Verkligen . 
Men kanske kassajobbet på Boans är värt att tänka på ? 
Du var fantastisk ! 
Hon är snäll , och han har ett ego stort som Moskva . 
Kanske . Men vi var ett bra team . 
Ja , det var vi . 
Jag måste be om en tjänst . 
- Vad som helst . - Kom ! 
Jag har ett problem . 
- Nu ! 
- Jag behöver en läkare . 
- Känner du någon ? - Det är klart . 
Men om du är sjuk , - borde Yvgeni veta ... - Jag är inte sjuk . 
Jag tror att jag är gravid . 
" Allt bra " , som ni australier säger ? 
Jadå , allt bra . 
Var har du varit ? 
Dansövning . Jag väntade på dig . 
Är du arg på mig ? 
Det var den tredje som du missade . 
Jag bara glömde . 
Förlåt . 
- Så du är inte ... 
- Arg ? Nej . 
Bra . 
Men du kysste min syster . 
Jag såg dig . Min lillasyster . 
Du skulle vara min vän . Eller hur ? Min medpilot . 
Vi och månen . 
Och du kysste min syster . 
Det hände bara en gång . 
- Jag är ledsen . 
- Två gånger . 
Jag såg er på taket . 
Jag försökte hjälpa henne . 
En gång , två gånger , 20 . Det kvittar . 
Hon är min lillasyster . 
Och du skulle vara min vän . 
Jag är din vän . 
- Tilly , det är jag . 
- Jaha . 
Det var bara ett dumt ögonblick , okej ? 
Och jag är ledsen . 
Jag trodde att du hade bättre smak gällande flickor . 
Jag har jättebra smak gällande danspartner ... Dansen ? Vem bryr sig om den jävla dansen ! 
- Jag trodde du ville dansa . 
- Jono , Mia dog nästan i krocken ... - Det är okej . - ... med min bäste vän . 
- Vi har löst det hela . - Nej . Det är inte okej . 
Mia är galen , mamma och pappa har tappat vettet , och någonstans där uppe är Skylab på väg ner . 
- Det är okej , Tilly . 
- Nej , det är det inte . 
Jag skrev till alla de där astronauterna , och ingen skrev tillbaka . 
- Astronauter ? De är upptagna . - Nej , det är de inte , Jono ! 
Ingen flyger till rymden längre . 
Ingen . 
Kom igen . 
NYHETER IKVÄLL Arbetare i Sydney protesterar mot fackföreningsgripanden . Beasley är ur form vilket pekar på mål till South Freemantle under veckoslutet , och miss Universum träffar miss Gerro ' . Tävlingen reser norrut . 
Godkväll , Perth . 
De sänder alltså inte historien . 
Bara Beasleys mål och miss Gerro . 
Inte lika viktigt som Bettys död . 
Det förtjänar en drink . 
Skandalen är begravd i arkiven . 
Jag slår vad om att det finns mer . 
Den lilla jäveln planerar något . 
Jag bara vet det . 
Pronto , tonto ! 
Skit . 
Vad fan var det där idag ? 
Nå ? 
Det var jag som fick sparken av min bror . 
- Jösses , Tony . 
- Förlåt . 
- Han avbröt dig och ... - Nej ! - ... jag tappade behärskningen . 
- Det gjorde du när han skymfade dig . 
Jag kvävdes av testosteronet i rummet . 
Och förresten - behöver ingen tala i mitt ställe . 
- Det stämmer . 
Hon klandrar mig jämt . 
Pappa . 
Det kunde ha varit en början på något nytt . Du och Mick . 
Det var det inte . Det var slutet . 
Men på plussidan ... Lillebror ger bra avgångsvederlag . 
Jag tog med Mia ut med den här . 
Hon älskade det . 
Oroa dig inte , imorgon ska vi surfa . 
Kom igen . 
Pappa . 
Den här sången påminner mig alltid om dig . 
Jag älskar den ! 
- Bara lyssna . 
Du är en starman . 
Det är du verkligen . 
Lovar du att aldrig släppa dina drömmar ? Då släpper jag inte mina , okej ? 
Okej . Men ... jag är en starwoman . 
Vad fan ? Vad ? 
- Vad vill du ? 
- Jag vill ge dig 1000 dollar så att du ger dem till din kompis , " Chicken " . 
- Chook ? 
- Chook . Chicken . 
Vänta lite . 
Du är pappan till den där tjejen . 
- Mia . 
- Ja . 
Hon krockade Chooks bil med den där asiatiske killen . 
Han är vietnames . 
Du är en av jävlarna som gör det svårt för våra familjer , va ? 
- Du , kompis ... - Va ? 
Här är pengarna till bilen . 
Säg till " Chicken " att ni kommer att lämna min dotter ifred . 
Och Jono . 
Och alla våra familjer . 
- Är det uppfattat ? 
- Chook . 
Skitstövel . 
Min bräda ! 
Jag åker först . 
Morfar ! 
Stig upp ! 
Morfar , snälla ! 
Snälla , någon hjälp ! 
Snälla ! 
PRODUCENTERNA TACKAR RESPEKTFULLT ABORIGINERNA OCH FOLKET PÅ TORRES STRAIT-ÖARNA DE SOM ENLIGT TRADITION ÄGER MARKEN OCH HAVET DÄR DETTA PROGRAM SPELATS IN , SAMT DERAS FORNA OCH NUTIDA ÄLDSTE . 
