Ta för er ! Hugg in ! 
Det är inte varje dag en mans dotter återvänder från de döda . 
Jag undrade varför alla tittade . 
I dag blev jag rånad av stråtrövare . 
Ringen på ditt finger . Du kanske måste donera den . 
En av dem slog mig . 
- Vem är du ? 
- Billy Blind . 
- Vad menar du med att du är på min sida ? 
- Jag skyddar dig . 
Jag är oåtkomlig . 
Charles Devereux , madam . Snobb . Bon viveur . Du är Isambard Tulley . 
Det hoppas jag inte . Han har en belöning på 20 pund . 
Pappa är död . 
Jag jagade ut honom ur stan i mörkret . Sen dödade jag honom . 
De försöker mörklägga det . Jag vill ha allt nu . 
Vad står mellan dig och din egendom ? 
Ska jag döda min egen far ? 
- Hon dödade honom ! 
- Nej , det gjorde jag inte ! 
Efter henne ! George , Roxy , vi sticker ! 
Vad händer ? 
Vart ska vi ? 
Jag berättar när vi är framme . 
Herregud , pappa . 
Hur kan du vara så arg på mig ? 
Det är alltid tumult i familjen när man gifter bort den äldsta dottern och nu måste stackars jag lida . 
Din mamma och jag har varit för fästa vid dig . - Pappa . 
- Om du inte får - mr Ledger som din älskare ... - Älskare ? 
Har han nånsin ens gett mig en försmäktande blick , skrivit en sonett eller kastat sig vid mina fötter ? 
- Varför gifta mig med honom ? - Han är en make som din far och mor tillhandahåller . 
Är de inte rätt personer att göra sig av med dig ? 
Göra sig av med mig ? 
Pappa , ditt huvud är så fullt av handel , att du skulle göra dig av med din dotter som en handelsvara . 
Mitt hjärta är min egen egendom och står bara till mitt förfogande . 
Hennes fräckhet förvånar mig . Din respektlösa slinka ! 
Inte respektlös alls , pappa ! Men sanningen är att mitt hjärta ... Så där . Nu är det sagt . 
Ser ni vilken situation jag är i ? 
Ingen bryr sig . Nonsens , jag tycker det är generöst av dem att dela sin smutsiga byk med oss . 
Du , sir , är full . 
Det är en väldigt ... Ja , det är jag . 
Herregud , pappa ! Vi har ökat farten ! 
Vi har lämnat huvudvägen . 
- Det är inte vägen till London ! - Spännande ! Vad händer ? 
Stanna maskinen ! 
Vad händer ? 
Herregud , pappa , vi har stannat . 
Ge mig den . 
Klä av dig nu . - Va ? - Kom igen . 
Du skulle inte hjälpa i slumpmässiga våldshandlingar , Billy Blind . 
Om någon riktar en pistol mot dig har jag skyldigheter . 
Det är bra att veta . Vänta . 
- Vilka skyldigheter ? 
- Jag vet inte . 
Var kom dessa skyldigheter ifrån ? - Nu ! - Det är en bra fråga . 
- Och svaret är ? - Knepigt . 
Jag måste anta att ditt liv är viktigt , eftersom jag ska skydda det . 
Men varför ? Varför ? Och fortsätt . 
Och vem bestämmer sånt ? 
- Du måste passa in på beskrivningen . 
- Som sagt , jag vet inte mer än du . - Kom igen . 
Skynda dig . 
- Ja , men du måste kunna ... 
- Vi ska inte ifrågasätta . 
Vi ska bara gå vidare . Ja , men ... 
Pappa , gör nåt . 
Billy ! Jag vill se hud . Kom igen , allt . Låt mig se det . Ut med dig då . 
- Ut med dig . 
- Jag sitter inte vid dörren . 
Jag är inte den enda vid dörren . 
Jag måste be om att bli ursäktad . 
Två saker , sir . 
Ett , vi vet inte vad som finns där ute . 
Och , B ... Jag är lite vek . 
Jag råder er att gå ut . - Av vem ? - Varför ? Upp med händerna . 
Hur står det till ? 
Lady Wilmot , överste Standring är här med en annan herre . Ja . Ta in dem hit . Säg åt min bror att komma ner . 
Jag vill inte behöva be två gånger . 
Thomas . 
Lämna mig ifred . 
Låt mig vara ! 
Blancheford . 
Lord Standring . Har du väntat länge ? Förlåt . 
Din syster har berättat att din förlust tar hårt på dig . 
Det måste ha varit en brutal attack . 
Jag beklagar sorgen , Ers nåd . 
- Det här är kapten Jarrold . 
- Hur står det till ? 
Om nån kan hitta din fars mördare är det Jarrold . 
Den här tiden i morgon har vi ögon i varje stad i England , lord Blancheford . 
Jaså ? 
Hur då ? 
Ni måste erbjuda en stor belöning . 
Vi annonserar i alla tidningar med en så detaljerad beskrivning av Nell Jackson som du kan ge och eventuella medbrottslingar . 
Vi får nyheter inom en vecka . 
Inom en månad kommer hon att hängas från schavotten . 
Att hitta henne är en sak . Att hålla fast henne är kanske nåt annat . 
Thomas har rätt , kapten Jarrold . 
Vi behöver mer kraft än du kan föreställa dig . 
Hon slåss tydligen som en demon . Och med tio mäns styrka . 
Hon är onaturlig . 
Jag ser fram emot det . 
Jag kan räkna löven från träden . Jag kan se enskilda föremål . Jag gillar inte att rota i andras saker . 
Jag gillar inte att sno andras saker . 
Jag gillar inte att vara i en position där jag måste sno andras saker . 
Ost . Vem vill ha ost ? 
- Kan jag få lite ost ? - Ja . 
Självklart , den är vår nu . 
Och jag bad dem om ursäkt . 
Jag sa att jag var i en svår sits som inte var mitt fel , och att jag har munnar att mätta . Jag omfördelade en del av förmögenheten . 
Vad sa de ? 
Du kommer att hängas . 
Inte mycket . 
Jag tänkte ändå inte dö i sängen . 
- Borde du inte ... - Ja , miss ? 
Binda fast oss ? Så att vi inte kan fly , sir . 
Jag har inget rep . Du får låtsas . 
Slösa inte dina sorger på dem , Roxy . 
De har mer saker än de behöver . 
Vet du vad som är vulgärt ? 
Varför behöver en man tio par byxor , medan en annan , en meter bort , måste gå nerför gatan med skinkorna hängande utanför byxorna ? 
Om världen var en bättre och rättvisare plats , skulle det här inte hända . 
- Jag vet . 
Jag vet det . - Jag vill åka hem . 
Jag har funderat på vad jag ska göra . 
Ingen av er har gjort nåt fel , - så i en god värld ... - Jag har det . 
Jag tog den här krabaten från lorden . 
Det är en enkelresa till det trebenta stoet , om det fanns någon . 
Det inte som det du gjorde , inte gjorde , men jag säger det bara . Jag hängs , precis som du , om de får tag på mig . 
Jag pratade med de här två , så jag tar itu med dig om en minut . 
Stick . 
I en god värld , skulle en rådman lyssna på sanningen . Men i den verkliga världen händer det inte . 
Så nu har jag mat i strupen , och jag kan tänka klart . 
Det vi borde göra ... är att åka västerut via småstigarna och de mindre vältrampade spåren , så släpper jag av er två hos farbror Jack i Abingdon . 
Är farbror Jack en riktig person ? Ja , självklart . Han är pappas lillebror . 
Du då , Nell ? 
Vad ska du göra ? 
När ryktet sprids om det här senaste rånet , tror de att vi är på Norra vägen . 
Så om vi åker västerut får vi ett försprång . 
Och när jag har släppt av er i Abingdon sticker jag till Bristol , smyger ombord en skuta - och seglar till Amerika . - Amerika ? 
Vad ? Ja . 
När jag har gjort mig hemmastadd och blivit något , skickar jag efter er . 
- Han då ? - Vem ? 
Ja , självklart . Ge mig en minut . 
Jag behöver prata med dig , här borta . 
Skynda dig . 
Vad är det , chefen ? 
Jag är inte din chef . 
Du måste ta tillbaka hästen . 
Skyll på mig . 
Säg att jag kidnappade dig , men sen lyckades du smita ifrån mig , okej ? 
Det här är inte din röra . Det är min . 
Men du måste tillbaka , så jag inte behöver oroa mig för dig och allt . 
Jag vill inte tillbaka . Jag skulle få stryk av pajasen Thomas . Okej . 
Åk inte tillbaka . Åk vart du vill . Men jag lämnar ungarna med tak över huvudet . Ingen kommer att se röken av mig . 
- Inklusive dig . - Varför ? 
Det är så det är . 
Vart ska du ? 
Ta för dig . Ta några fina , varma plagg . Ta ett par . 
- Kan jag inte bara hänga med dig ? - Nej . 
Kan jag inte vara till nytta för dig ? 
- Nej . - Om du hade låtit mig följa med och ta vagnen i morse hade du sett hur användbar jag kan vara . 
Ja . Jag tillhör ingen duo . 
Jag försökte med kapten Jackson och jag lärde mig är att det är var man för sig själv . 
Men se , du är fri . 
Världen ligger för dina fötter . Som du med svärd kan öppna , va ? 
Ja , greppa den . 
Världen är stor . Det finns mycket att se och göra . Du får sätta fart . 
Sätt fart . 
- Gratulationer är på sin plats . 
Du fick som du ville . Marken , egendomen , titeln . 
Du är en rik man , Blancheford . Och en så enkel lösning . 
En som fanns där hela tiden , bara väntade på att bli tagen . Snälla . 
Det låter som om du kom undan med det , eftersom alla skyller på den här kvinnan , Nelly Jackson . - Ja . Bra gjort . - Jag ... 
Lappen bad mig söka upp dig . 
- När är begravningen ? - I morgon . 
Jag kommer . 
Du kände inte min far . 
Begravningar är inte för de döda , Thomas . 
Jag ska stötta dig och din syster 
- i er mörka timme . 
- Du känner inte min syster . 
Jag såg henne vid hovet för ett antal år sedan innan hon gifte sig med lord Wilmot . 
Stackars karl . Stackars flicka . Hon sörjer fortfarande sin make . Nu har hon förlorat sin far . 
Begravningsprocessionen lämnar huset klockan sju . 
Men du behöver inte ... Jag vill . 
Du förstår , folk som du är sällsynta , Thomas . 
Jag visste inte om du var kapabel . 
Jag var inte säker på att du inte var en bortskämd liten pojke . Men nu är jag nyfiken . 
Jag känner ett visst ansvar för det som hände . Men jag undrar vad mer du är kapabel till ? 
Jag undrar om du inte är skapt för stora saker . 
Vad för saker ? 
Det kommer en tid för det . 
Jag ville bara veta när begravningen var och jag ville träffa dig . 
Jag har saker att göra . Vi ses i kyrkan . 
Benning följer dig ut . 
Han måste sätta sin prägel på världen och Rasselas kan väl inte göra det om han tramsar runt med oss ? Nej . 
Han måste göra vad han kan med sitt liv medan han har chansen . 
- Men jag gillade honom . 
- Jag gillade honom . 
Jag gillade honom . 
Ja , men jag menar ... Jag gillade honom . 
Ja , men den sortens sörja är en lyx vi inte har råd med just nu . Det vore en olägenhet . Och risken finns med sånt här , att båda inte känner likadant . Jag vill inte se dig förkrossad . Han gillade mig . Han sa det . 
Gjorde han ? 
Så olämpligt . Han borde ha hållit det för sig själv . 
Jag misstänker att han är åtta , - tio år äldre än du . - Tre . 
- Tre år äldre än jag , det är allt . - Och ... 
- Du är inte min mamma . - Och ... 
Nej , och det vill jag inte vara . Jag har aldrig sett nån vara så snabb . 
Så när har ni haft alla dessa djupa samtal då ? 
Här och där och längs vägen . 
Och hans far var , tja , är kungen av Benin . 
Verkligen ? 
Ja , det är troligt . 
Det säger han säkert till alla dumma 16-åringar med lite ludd mellan öronen . 
Varför berättade han vad han hade hört - om vad som pågick ? - Jag vet inte . 
Varför skulle han riskera livet om han inte brydde sig om folk ? 
Han hade sett mig i byn och tyckte att jag var ... 
En engelsk ros . 
Vad är det då ? Har ni kyssts ? - Nej . - Visst . - Vem har kyssts ? - Vi har pratat . - Hon och Rasselas . - Ingen . Ingen har gjort mer än att lyssna på livshistorier . - Jag vet inte . 
- Det var det jag sa . Han köptes i Londons hamn . 
Tre år gammal för 15 pund , åtta shilling och sex pence av lord Blancheford . Han tog mig tillbaka till Tottenham på sin häst . 
Det var åska och blixtar . Lord Blancheford höll mig varm under sin mantel . Jag tvättades och kläddes och gavs till Sofia och grisen Thomas som leksak . 
De hade just förlorat sin mor . Lord Blancheford ville muntra upp dem . 
Han fick mat ... kläder och blev klappad och behandlad som en i familjen , tills en dag ... När Rasselas var nio eller elva ... Thomas skickades till Eton eller nåt sånt , och jag sattes i arbete på gården . 
Miss Sofia och Rasselas grät och grät , men ... Det var då allt förändrades , och ... Pengarna eller livet ! 
- Ut ! - George , kom . Vad händer ? 
- Ut , sa jag ! 
- Nell , vad händer ? 
Det är tomt , guvernören . 
Det är bara en massa kläder . Vänta lite . 
- Jag känner dig . 
- Det gör du . Varför inte plåga nån annan innan jag benar ditt hår som sist ? 
Och vilka är de här två skönheterna ? 
Det är den där karln , Nelly . 
Den där snobben från London . 
Vad försöker den stackaren säga ? 
Det är vi , mr Devereux . 
Varför är du klädd som en stråtrövare ? 
Vad hon försöker säga är , jag träffade en kille i London som är otroligt lik dig . 
Man skulle kunna tro att ni var tvillingar . 
Han hade till och med ett ärr , som jag kunde svära på att jag gett dig , honom , själv . 
- Märkligt . 
- Hur kom du över den här vackra vagnen - och de här fyra hästarna ? - Jag fick låna dem . 
Vet du vad jag tror ? 
Jag tror att du är Nelly Jackson . 
Nelly Jackson , som har en belöning på 20 pund på sitt huvud för mord . 
Det tog mig 18 månader att få en belöning på 20 pund . Den här gör det på en natt ! Hela London vet om det . 
I morgon kommer det att vara upp , ner och i sidled över hela landet . 
- 20 pund ? 
- Vad sägs om det ? Vi tar den här hästen , de fyra hästarna och vagnen och de här två slamporna , och lämnar in den snacksaliga och får de 20 punden . 
Har ni inte lärt er något från förra gången jag spöade upp er ? 
Iväg . 
Han är ny . 
Det är logiskt . 
Kom igen då . 
- Släpp pistolen . - Rasselas ! 
Vad ska jag göra med den här ? 
- Vad gör du här ? 
- Jag räddade dig . Förlåt . 
Räddade du mig ? 
Vadå " räddade mig " ? 
Och Roxy och George . 
Följde du efter oss ? 
Så jag tänkte gå min egen väg , som du föreslog . 
Men jag ska vara ärlig , chefen . Jag kände mig ledsen . Sen kände jag mig ensam . Sen kom jag hit och oroade mig för er tre , och ... Vad ska jag göra med honom ? 
Jag vet inte . 
Det beror på vilken smörja som kommer ut ur hans rövhål härnäst . 
Jag kunde inte erkänna att jag var Charles Devereux inför akademikerna , eller hur ? 
Vad hände sen ? 
Gick du tillbaka och dödade avskummet som mördade din pappa ? 
Nej , det gjorde jag inte . 
Det är vad alla tror . Jag har en idé . Du kommer att åka fast . Jag vet inte din plan , men eftersom vi står här mitt på dagen och diskuterar det här , så antar jag att den är dålig . 
Jag hoppas du inte lämnar småttingarna hos en favoritfarbror , Nell ? 
Inte den gamla godingen , väl ? 
Även om jag gjorde det , vilket jag inte gör ... 
Där letar de först . 
Om du har en syssling som du aldrig har sett , som bor i Kent , står de utanför hans hus i morgon . 20 pund är mycket damm . 
Vill du höra min idé ? 
- Det kan jag göra . 
- Vi borde slå ihop oss . - Nej . 
- Jag kan hjälpa dig . 
Det tvivlar jag på . 
Som jag sa , vid den här tiden i morgon kommer alla nyhetsblad i landet att trycka din beskrivning , och inte bara din , hennes och hennes och hans . 
Det finns ingenstans ni kan gömma er . 
Så vad gör du ? 
Vart åker ni när det inte finns någonstans att ta vägen ? 
Fick du nån kosing när du lånade den här benströaren ? 
Några pund , kanske . 
Vi låtsas vara lord och lady si och så och hyr bra rum på ett fint hotell i en likgiltig stad i några dagar . 
Du har kläderna . Låt oss använda dem . Vad pratar du om ? 
Jag pratar om att gömma oss helt öppet , Nelly Jackson . 
Det innebär att inte gömma sig alls . Man förändrar bara den man verkar vara . 
Vi då ? 
Hennes nåd måste ha en kammarjungfru . 
Hennes nåd kanske reser med sin excentriska lilla kusin . Och lord Den-och-Den måste ha en bra lakej . Ja , eller så kan du vara min lakej . 
Tänk bara . Varm mat . Varma sängar , rena kläder , tak över huvudet . 
Varför ? 
Varför gör du det ? Vad får du ut av det ? 
Jag gillar äventyr . 
Alla tittar på mig . 
Nej , det gör de inte . 
Jag är uppståndelsen och livet , säger Herren . 
Den som tror på mig , skall leva om han än dör . 
Och den som lever och tror på mig ... skall aldrig dö . 
Jag vet att min förlossare lever och att han till slut skall stå fram över jorden . 
Inga maskar förgör denna kropp . Thomas . 
Genom mitt kött skall jag se Gud . 
Fortsätt bara . 
Som jag skall se med egna ögon och mina skall jag skåda . 
Vi hade inget med oss till världen och det är säkert att vi inte kan ta med oss något ut ur den . 
Välsignat vare Herrens namn . 
Amen . 
Amen . 
Lord och Lady Shankley . 
Ja , det är vi . 
Anmärkningsvärt anskrämlig . 
- Är det en kvinna ? 
- Självklart är det det . 
Bathsheba . Barn ska synas men inte höras . 
Får ni inte kalla kårar av hennes uppsyn ? 
Tvärtom , det är det andra som gör mig nervös . 
Ser du hur ett av hans ögon är mindre än det andra ? 
Ja , ma ' am . Ganska groteskt . 
Jag ser inte det . Men hon är ganska sjaskig . 
Luktar han till vänster illa ? 
Ja . 
Det är första gången någon vill ha henne . 
Mycket bra . Jag vill slå honom på käften . 
Tänk att vara stråtrövare . 
Tycker du att hon är vacker ? - En hagga . - Dumma hatt . 
Ser ut som en vessla . 
Ser hans näsa ut som en hunds snorre ? 
Håller du med ? 
Vad tycker du ? 
EFTERLYST AV DROTTNINGEN . ISAMBARD TULLEY , BELÖNING PÅ 20 PUND EFTERLYST AV DROTTNINGEN . Båda är lika fina , sir . Våra rum ? 
Den här vägen , lord Shankley . 
Bagaget , Jacques ! 
Framåt ! 
Jacques . 
Ursäkta mig , mina herrar . 
Ursäkta , min gode man . Var hittar jag frun i huset ? 
Den här vägen , sir . 
Ja . 
Lady Wilmot . 
- Jag beklagar sorgen . - Har vi träffats ? 
Jag är Robert Hennessey . Greve av Poynton . 
Jag visste inte att min far kände någon i riksrådet . 
Det gjorde han inte . Inte mig i alla fall . 
Din far skickade din bror till London till din farbror James Ogilvy , din avlidna mors ... Min mors bror , ja . Ja , för att se om han kunde ... göra något med Thomas . 
Jag hade en bortkastad ungdom själv . Ogilvy trodde väl att jag kunde bli nån sorts guide , eller mentor åt Thomas . 
Det visste jag inte . Så vänligt av dig . 
Jag avbröt dig . 
Jag försöker bekanta mig med egendomsfrågor . 
Thomas gör det inte , men jag låter det inte gå till spillo . 
Om jag kan göra något för att vara till nytta , så fråga bara . 
Den enda nyttan någon kan göra är att ställa de depraverade icke-väsen inför rätta som mördade min far . 
Nell Jackson ? 
Frun . Mr Jarrold är här . 
Han säger att han vet att det är fel tillfälle ... 
Visa in honom . 
Jag har anlitat Jarrold för att spåra upp henne . 
Han är tydligen väldigt bra , men jag tror att det krävs mer än vanliga dödliga för att fånga henne . 
Har Thomas berättat ? 
Hon slåss som om ... hon är besatt av en demon . 
Och du såg det ? Såg du henne döda din far ? 
Ja . Hon sköt honom . Mitt framför oss . 
Kocken och några av männen sprang in när Thomas skrek , och ... Det var otroligt . Hon stoppade kulor med sina bara händer . 
Har du ... hört talas om sånt ? 
Det finns fler saker i världen än de flesta kan föreställa sig . 
- Verkligen ? 
- Ja . 
Det låter som att Nell Jackson kan ha , vare sig hon vet det eller inte , fått tillgång till en ande . Ett väsen . 
Och om hon har det , måste lika bekämpas med lika , för som du har sett , kan ingen dödlig röra henne . 
Kan du hjälpa oss ? 
Kanske . 
- Lady Wilmot . 
- Ska jag ... Stanna , är du snäll . 
Jag fattar mig kort . 
I morse hörde vi om en vagn som stoppats av en kvinna söder om Potters Bar . 
Att döma av hennes utseende och sättet hon uppförde sig på , så var det hon . 
Det kommer fler observationer . Och då kommer nätet att dras åt . 
Var hon ensam ? 
Vakten och föraren var tungt beväpnade . 
Båda var före detta soldater . 
Sätt in fler annonser i fler nyhetssidor . Och höj belöningen till 40 pund . 
Mycket bra . 
Bra , det är mycket bra . 
Lady Shankley , titta . 
Ja . 
Jag kunde ha varit i Bristol nu . På ett skepp . 
Saken är den , att jag inte borde känna mig tvungen att fly . 
En rådman borde lyssna på sanningen . 
Det kommer inte att hända . 
Lagen är skapad av snobbar för snobbar . - Sanningen är irrelevant ... - Visst . Eller det de vill att den är . 
- Det borde inte vara så . 
- Men det är så de tänker . 
Du hittar ingen annorlunda . 
Varför lever du så här om du är rik ? 
Du antar att jag har ett val . Jag är pank . 
Nej , det är sant . 
Farsan gillade spelborden för mycket . Lämnade mig nästan inget . 
Bara titeln och min adress i Mayfair , som jag är väldigt förtjust i . Förutom att det är fullt av hyresgäster . Jag har bara två rum på vinden . 
Men än sen ? 
Det är en adress i Mayfair ! 
Det är allt som räknas . 
Om folk kan ha förtroende för dig , för den du säger att du är , får det dem att känna sig bekväma . Då kan du komma undan med nästan vad som helst . 
Lysande . 
Nelly trodde mig inte när jag sa att din pappa var kungen av Benin . 
Oftast tror jag det knappt själv . 
- Men du känner dig lurad ? - Ja . 
Och mitt namn också . 
Rasselas är inte mitt namn . Lord Blancheford gav mig det . 
Mitt riktiga namn är borta , som min familj . 
Har du aldrig velat åka tillbaka och hitta dem ? 
Det skulle jag , mer än något annat . Men hur ? 
Jag vet inte var jag skulle börja även om jag sparade till resan . Och med allt som har hänt , om jag går i närheten av hamnen , sätter någon bojor på mig , och jag kan skickas till kolonierna . 
Det måste finnas ett sätt . 
Jacques ? 
Ett meddelande till din guvernör . 
Ett , två ... Gå då . 
Tack , lakej . 
Jag är inte din lakej , din ficktjuv . 
Jag låtsas vara din lakej . 
Det är en inbjudan till lord och lady Shankley att spela kort i morgon eftermiddag på Widdicombe Manor - med lord och lady Springbourne . - Vilka är det ? Vi träffade dem i kyrkan i går . Vi pratade med honom . 
Jag gjorde det . 
Jag sa att vi var på genomresa på väg till London och de har gjort det hövliga och bjudit in oss på te och kortspel . 
Du måste skriva tillbaka och säga att vi inte kan gå . Varför ? 
När jag öppnar kakhålet kommer de nog att märka att jag inte kan skilja ena ändan av gaffeln från den andra . Nelly , du är en sån besvikelse . Vi kan skinna honom vid spelbordet . - Jag kan inte . 
- Jag kan . 
Vi kommer att tjäna storkovan . 
Du var förvånansvärt övertygande som lady Shankley när vi kom , Nelly . 
George har rätt . Du har en naturlig ... - någonting med dig . - Jag tog med den här också . Ifall det står något om dig i den . 
Se det så här . Ju mer du övar på att låtsas vara nån annan , desto bättre blir du . 
Dessutom , Nelly , lord Springbourne , kan vara rådman . 
Du kan se vad han är för typ , om han verkar lyssna bra ... - När väntar de oss ? - Klockan fyra . 
Lyssna på det här . 
" Skurken som rånade och stal en vagn utanför Potters Bar för tre dagar sen , tros vara samma Nelly Jackson som begick mordet på lord Blancheford . " 
Varför kallas jag Nelly ? 
" I så fall kan man anta att odjuret ... " Är det du ? - Ja . - " ... är på väg norrut . " De har fel . Om alla tror att vi är på väg norrut , kan vi klara oss här i Slough i en vecka . 
" Belöningen för information som leder till gripandet av Jackson har höjts till 40 pund . " 
Poynton . Poynton ! 
Har du hållit dig uppdaterad om Nell Jackson ? 
Det är nåt övernaturligt över henne . 
Jaså ? 
Jag trodde att det var ditt expertområde . 
Jag undrade om hon kunde vara till nytta för saken . 
Jag hoppas att det är upp till mig att avgöra . 
Ja , självklart . 
Min chef tyckte det var nåt skumt med dem . Så fort de dök upp , tja , så fort hennes nåd öppnar munnen , och försöker prata som en sprätt . 
De sa att de var från Thunderbridge Hall i Totnes , men mrs Blewitt , som jobbar i köket , kommer därifrån och har aldrig hört talas om Thunderbridge Hall . Inte om lord och lady Shankley heller . 
Jag vet inte vem lord Shankley är , men beskrivningen av de fyra andra passar perfekt , inklusive rymlingen Rasselas . 
Pojken såg en lapp där de bjöds in på te i eftermiddag hemma hos lord Springbourne . 
Vad väntar du på ? 
Ge dig av nu om du vill fånga dem där . 
Kom igen . 
Får jag en del av belöningen ? 
Hur kan jag kontakta din vän , greven av Poynton ? 
Varför ? 
Det måste se ut som om vi gör allt vi kan för att hitta Nell Jackson . På grund av den idiotiska röran du försatte oss i . - Ja , men ... - Om du hängs för mord , går godset till vår kusin i Northumberland . 
Han flyttar in med sin familj och jag blir beroende av honom för varje smula . 
Så var stark . 
Bestämd . 
För min skull . Jag kan bara hjälpa dig om du hjälper mig . 
Mr Jarrold ? 
Jag ska skriva en lapp till greven av Poynton . Men sen vill jag följa dig och dina män till Slough . 
Gör dig redo . 
Kom igen . 
Kom igen . 
- Hur länge har vi varit gifta ? - Hur länge har vi varit gifta ? 
- Sex månader . 
- Sex månader , tre veckor , tre dagar . 
Detaljerna är viktiga . - Vad är min favoritmat ? 
- Ål i gelé ? Vaniljsås ? 
Kanderat äpple , kvitten , plommon och kalebass . Och kryddiga läckerheter från silkeslena Samarkand . 
Ska jag komma ihåg allt det ? 
Jag litar på dig , lady Shankley . 
Från början , min kära . 
Ett brev till er , sir . 
Det är inte så illa att vara på rymmen . 
Jag saknar inte den varma , svettiga tvätten hela dagen . 
Jag undrar hur Nelly började slåss så där ? 
Tror du att kapten Jackson tar hand om henne från andra sidan ? 
Det är något . 
Jag såg det . 
Hur då ? 
Jag vet inte . 
- Hur ser det ut ? - Det är som ... en aura . 
- Jag vet inte . 
- Vad har du sett ? Och den är bra . Den känns bra . 
Jag vet inte om kapten Jackson var bra . 
Är inte det lady Wilmot ? 
De vet att vi är här . Hur då ? De stannar inte . 
De vet att Nell är på Widdicombe Manor ! 
Hur då ? De är för många . 
Vad ska vi göra ? 
Fickdykare . 
- Vad är min favoritfärg ? 
- Typ , brun , lite dyngfärgad ? Akvamarin . 
Det här är ett misstag , Nelly Jackson . 
Upp med hakan . Se inte ner . Se folk i ögonen och le . 
Jag är inte säker på detta . 
Nonsens . Om du tvekar , titta bara på mig som om du är kär , så kommer jag på nåt . Jag säger dig , Nelly . Något konstigt kommer hitåt . 
God eftermiddag , och vilken strålande eftermiddag det är . 
