Seongmin . 
Titta , det är havet . 
Där , där . 
- Samsik . 
- Ja ? 
Ser du skeppet där borta ? 
- Ja , herrn . - Vad tror du driver ett så stort skepp ? 
Olja . Det är olja . 
Att sälja olja är det enda sättet att bli riktigt rik . 
Uncle Samsik 
Uncle Samsik 
Den avlidne Den 6 mars 1960 Seoul , Sydkorea Demokratiska partiet 
- Han kommer . - Han är här . 
- Här kommer han ! - Herrn ! 
Har ledamot Kang bett om ursäkt ? 
Ska du anmäla honom till etikkommittén ? 
Vad gjorde du i Nationalförsamlingen ? 
Kände du redan till om deras plan för lagförslaget ? 
- Vi går . 
- Kom nu . 
Vi fördömer starkt att lagförslaget antogs så skyndsamt och begär en officiell ursäkt från ledamot Kang och Liberala partiet . Annars måste vi klaga hos etikkommittén . Jag ber om ursäkt . 
Officiellt . 
Då röstar vi om lagförslaget igen . 
Ändringen för lokalt självstyre är redan godkänd . 
Men genomförandet var olagligt ! 
Det räcker . 
Då begär jag att du officiellt ber om ursäkt till ordförande Kim San . Samt publicerar en ursäkt i Liberala partiets nyhetsbrev och nyhetstidningar . 
Det är onödigt . 
Jag godtar hans ursäkt . 
Va ? 
- Du kan inte släta över saker . 
- Jo , ibland . 
Det räcker . 
Varför gjorde du så ? 
Det är okej . 
- Jag hör av mig . - Vänta . Vänta . 
Du skulle vara snäll mot honom . 
Jag menar ... Han slog nån i Nationalförsamlingen . 
Hur skulle jag annars se ut ? 
Kollade du listan jag skickade ? 
Ja , men ... 
Låt oss diskutera medlemmarna i Högsta rådet och de lokala ordförandena igen . 
Vi har redan en överenskommelse . 
Gör som jag säger . Och boka ett möte med Kang Seongmin . 
Jag övertalar mitt parti att inte gå till etikkommittén . 
Det var allt . 
Har du en minut ? 
Yeojin . 
Vad hände ? 
- Vad menar du ? 
- Är du journalist nu ? 
Jag studerade ju litteratur trots allt . 
Det här är obekvämt för oss båda . 
Det blir det inte om du håller dig i skinnet . 
Kom igen , Yeojin . 
Vi borde åka . 
Han har somnat . 
Vi väcker honom inte . 
Hans tillstånd var kritiskt i morse . 
Han klarar sig säkert . 
Kan jag leva upp till min far ? 
Ursäkta ? 
Ja , självklart . 
Jag är faktiskt rädd att jag ska förstöra min fars bedrifter . 
Jag hjälper dig . 
Han har varit förbundets mittpunkt länge . 
Allt löser sig med det parlamentariska systemet . 
Blir reformen av ? 
Självklart . 
Jag ska träffa ledamot Sun Wooseok . 
Varför vill du diskutera det ? 
Du har gått med på villkoren . 
Jag vill diskutera igen . 
Säg inte att du plötsligt har ändrat dig . 
Kom igen , var inte löjlig . 
Lista över kabinettsmedlemmar Valkretsarnas fördelning 
Det här är inte bra . 
Våra medlemmar har suttit över tre mandatperioder . 
Det spelar ingen roll . 
Ni har de viktiga rollerna medan vi har smulorna . 
Vi är över 100 personer . 
Högsta rådet måste delas lika . Vi utser tre ministrar och vice ministrar inom ekonomin . 
Tänk på att vi är överlägset fler än ni . 
Kan ni säkra fler än 100 platser ? 
Jag kan säkra trettio platser från Demokratiska partiet . 
Mitt svar är nej . 
Ärligt talat finns det folk som hyser misstankar mot dig . 
Vilka misstankar ? 
Jag menar ryktet om Sineuialliansen . 
Vem tror på det grundlösa ryktet ? 
Inte jag , så klart . 
Så vem gör det ? 
Ge oss deras namn . 
Om An Yosub misstänker honom , vänder Cheongwooföbundet honom ryggen . 
An Yosub klarar sig inte länge till . 
Jag såg honom på sjukhuset . 
Hans dagar är räknade . Och vad kan den där ungen , An Kichul , göra ? 
Vi har Cheongwooförbundet under kontroll . 
Vad håller du på med ? 
Vad i hela friden pågår ? 
Vill du dra dig ur ? Är det så ? 
Vad sa du till mig ? 
Varför gör du så här ? 
Var kommer detta ifrån ? 
Tror du att det är lätt att förena två partier ? 
Säg inte att du har ändrat dig . 
Jag vill förhandla lite till , okej ? 
De har alla suttit över tre mandatperioder ! 
Inget av det här är lätt ! 
Jag räknar med dig . 
Oroa dig inte , herrn . 
Han spelar bara svårfångad . 
Han ser ner på mig . Han tror att demokraterna vinner . 
Både Cheongwooförbundet och Liberala partiet vill överge mig . 
De jävlarna bryter sitt löfte för att jag är mesig . 
President Rhee vinner säkert . 
Tänk på hur Choi Minkyu är . 
Han skyr inga medel . 
Sun Wooseok backar när valet är över . 
Jag tror inte att presidenten vinner . 
Du , det går att vinna . 
Hur då ? 
Den avlidne Choo Intae . 
Ska vi använda en död person ? 
Vi använder honom eftersom han är död . 
Demokratiska partiet 
Kom in . 
- Ville du träffa mig ? - Ja . 
Jag har gått igenom utkastet till dina löften . Partimedlemmarna godkände det . 
Jag går händelserna i förväg , men båda partigrupperna jobbar på strukturen för nästa kabinett . Ledamot Sun föreslog ett ministerie för nationell rekonstruktion . 
Vad säger du ? 
Så istället för inrikesministeriet ... 
Du kan väl börja planera strukturen ? 
Jag la ett gott ord för dig . 
Vi pratar här . 
Jag vet att ditt mål är att implementera rekonstruktionsprojektet . 
- Tack så mycket . 
- Vem vet ? 
Du kanske till och med blir minister för nationell rekonstruktion . 
Det vore en dröm . 
Kan vi implementera det parlamentariska systemet ? 
Jag frågar farbror Samsik . 
Varför ska du diskutera det med honom ? 
Lita inte för mycket på honom . 
Han är en vältalig orm . 
Håll tyst runt honom . 
Ledamot Sun gav upp parlamentssystemet . Av goda skäl . 
Demokraternas popularitetssiffror var skyhöga . 
Höll du det hemligt för Samsik ? 
Nej . 
Varför inte ? 
Välkommen . 
- Ge oss lite whisky . 
- Okej . 
Den vanliga , herrn ? 
Visst , det låter bra . 
Ska bli . 
Du verkade populär på kampanjmötet . 
Kom igen . 
Väljarna stöttar vem som helst från vårt parti nu för tiden . 
Du borde ändå gå på fler möten . 
Du måste träna mer för att hänga med . 
Jag vet . Men tyvärr är sex min enda träning . 
Så du tränar bara två minuter i månaden ? 
Hallå . 
Eller en minut ? 
Det är bättre än inget . 
Man måste vara i form för att röra sig mellan två sidor . 
Vad är det med dig ? 
Vi pratar utanför . 
Vad gäller det ? 
Har Kang Seongmin sagt nåt ? 
- Vad sa du till Kim San ? 
- Va ? 
Försökte du locka honom med en ministerroll ? 
Så han har redan skvallrat ? 
Han berättade inte om dig . Han försökte bara övertala mig . 
Han sa att han inte bryr sig om positioner . 
Han vill hindra min förening med Kang Seongmin . 
Så oskyldig är han . Hur kan du locka en sån man ? 
Skäms på dig . 
Din ytlighet håller dig i utkanten . 
Jag försökte inte dra mig ur . 
Ska jag berätta för alla om föreningen med Kang Seongmin ? 
Förlåt . 
Försök inte övertala honom igen . 
Okej . Jag ska vara försiktig . 
Föreningen sker som överenskommet . 
Visst , jag förstår . 
Okej . 
Samsik var emot idén om ett ministerium . 
Så varför berättade du ? 
För att ni saknar hemligheter ? 
Varför berättade du allt ? 
- Bra jobbat i dag . 
Vad gör du här ? 
Har du en minut ? 
Vi måste prata . 
Jag borde ha undvikit Yoon Palbong och Innovationspartiet . 
San . Jag är glad över Cheongwooförbundet , men orolig över de senaste händelserna . 
Jag behöver din hjälp . 
Säg till farbror Samsik att jag inte klarar det . 
Jag pratar med honom så att han förstår . 
Oroa dig inte , okej ? 
Var har du varit ? 
Jag hade ett middagsmöte . 
- Du borde gå hem . 
- Okej . 
Du har jobbat hårt med lutfabriken . 
Det har jag . 
Tänker du kasta bort allt hårt arbete ? 
Nej , herrn . 
Vi vill väl ... att Kim San ska bli premiärminister ? 
Självklart . 
Det finns inget värre än halvfärdiga jobb . 
- Jag ... 
- Hindra inte din vän . 
Jag är livrädd . 
Ta dig samman , okej ? 
Vill du så gärna hindra minister Kim ? Vill du det ? 
För ett hederligt liv behövde du släppa din girighet . Men du ville ha både lutfabriken och Cheongwooförbundet . 
Man får bara tillfredsställa några begär . 
Ingen får alla . 
Det är givet . 
Så vad ska vi göra ? 
Du borde öka dina begär . 
Har du inga ambitioner ? 
Du planerade en statskupp hela tiden , va ? 
Det var därför du berättade allt för Samsik . 
Nej . 
Jag planerar en statskupp . 
Kapitalförsvaret , 3:e marinkårsregementet , 55:e Howitzerregementet , och en dödspatrull på 30 man från armén . 
Efter presidentvalet åker presidenten till sitt fritidshus . 
Om vi tar honom som gisslan , förklarar undantagstillstånd och blockerar vägarna till huvudstaden , finns det hopp . 
Jag kan inte låta vårt land hamna i fel händer igen . 
Jag planerade inte att genomföra en statskupp . 
Men det gjorde du . 
Om du misstrodde mig från början varför kom du till rum 806 på Hotell Banya ? 
Och varför bjöd du in mig ? 
Jag tycker att vi är kvitt . 
Hej , herrn . 
Tack för att du kom . 
Rachael Jeong från Albright . Trevligt att träffas . 
- Är general Choi här ? 
- Ja , där uppe . 
Den här vägen . 
Vi var båda tveksamma och frågade ut varandra , väl ? 
Precis . 
Planen lät genomförbar . 
Drick upp . 
Presidentens fritidshus vaktas vanligtvis av 20 personer . Den 122:a bataljonen kan ta sig dit inom en timme . 
- Vi måste hålla de borta . - Ja . 
Vi behöver logistikkommandots hjälp för att flytta trupper och utrustning snabbt och diskret . 
Vi börjar förbereda när datumet är satt . 
Planen verkade perfekt och lagom berättigad . 
Varför inledde du inte statskuppen direkt ? 
Den skulle ju ske . 
Om du var i min sits vad hade du gjort , överste ? 
Vi soldater har strategier baserade på resurser . 
Vi förlitar oss inte på antaganden om en möjlig vinst i valet eller införande av parlamentssystem . 
Så är soldater . 
Var inte du själv soldat ? 
Minns du den dagen ? 
Väldigt tydligt . 
Det var en hektisk dag . 
Det var min idé att etablera Albright . 
Jaså ? 
Min far uppmuntrade mig att prova nåt i Korea . 
Det var utmanande först , men jag gillar det . 
Skönt att höra . 
Det är min farbror . 
Farbror , senator Jeremy Albright . 
Han är utrikesminister . 
Han har varit till stor hjälp . 
Jag har träffat honom förut . 
Farbror Jeremy talade väl om dig . 
Gjorde han ? 
Ursäkta mig . 
General Choi har gått . 
Tack . 
Mötet är avslutat . 
Bra jobbat . 
Nu kan jag slappna av . 
Har du en cigarett ? 
Så minister Albright talade väl om mig ? 
Han sa att du var vår bästa alumn . 
Det sa alla andra också . 
När jag studerade i USA gjorde jag allt för att överträffa de framstående eleverna . 
Så alla sa till mig att jag kunde förändra Korea till det bättre och att det var min plikt mot mitt land . 
Men tänk att det skulle ta sån tid . 
Så det är det du är rädd för . 
Det är nog inte för sent . 
För dina idéer , dina åsikter och din vision om ett nytt Korea ... Det har öppnat mitt sinne . 
Jag tror faktiskt att du kan förändra allt . 
Jag ska vara ärlig . 
Jag har en bekännelse . 
Vadå ? 
Låt höra . 
Jag tog in general Choi . 
Va ? 
Och jag valde dig . 
Jag tror inte att Korea är redo för demokrati . 
Därför behövs en utmärkt ledare . 
Jag fick den drömmen när jag kom hit . 
Att fostra en bra ledare . 
En eminent ledare . 
Du har tur . 
Jag har inget val . 
Varför välja nån annan ? 
Välj mig , så följer familjen Albright med . 
Tack . 
Säg inte till farbror Samsik att du träffade general Jang . 
Vi får väl se . 
Verkade Choi Hanrim omedveten om allt ? 
Ja . 
Vill du ha bröd ? 
Jag vill ha vatten . 
Visst . 
Jag träffade precis ledamot Sun Wooseok . 
Det gör väl inget ? Nej . 
Ta inte åt dig av det han sa . 
Folk ger alla möjliga löften under val . 
De ska röra upp himmel och jord och lovar all möjlig makt . 
Jag gick inte på det . 
Har det hänt nåt bra ? 
Nej . Hur så ? 
Du verkar vara på bättre humör än vanligt . 
Jag tog några drinkar bara . 
Med vem ? 
Rachael . 
Bjöd hon ut dig på en drink ? 
Hon ville fördriva tid i väntan på general Jang . 
Hon måste gilla dig . 
Varför stöter du inte på henne ? 
Det vore betryggande att ha familjen Albright bakom dig . 
Låt oss prata affärer . 
Pak Jiwook kommer att anmälas i morgon . 
Jag förstår . 
Är vi klara ? 
Minister Kim . 
Jag är glad att se dig på så gott humör . 
Bjud mig på en drink , då . 
Visst , det ska jag . 
Jag ringer dig . 
Det fjärde presidentvalet , som äger rum den 15 mars , är runt hörnet . 
Båda kandidaterna har kampanjat nonstop för att få väljarnas stöd . 
Med Demokratiska partiets ökande popularitet , har partiet lagt fram ny ekonomisk politik för att skilja sig från nuvarande administration . 
Folk samlade i Jangchungdan applåderade demokraternas politik . 
Flera politiska kommentatorer sa att liberalerna behöver väljare på landsbygden för att president Rhee ska få sitta en period till . 
Rösta på nummer 1 
Rhee Seungmin som president Rhee Kihak som vice president 
Rösta på nummer ett ! 
- Nummer ett ! - Nummer ett ! 
När det lokala självstyret har ändrats utses personal till alla lokala regeringar . De kommer att samla in valsedlar från äldre , tidigare invånare och valskolkare för att säkra 40 % stöd före valet . 
Kom ihåg era tilldelade grupper och följ planen på valdagen , okej ? 
Vilken grupp ... 
Du är i min grupp . 
Hallå där ! 
Ni ska vara i grupper om tre ! 
Är det ett skämt för er ? 
Kom hit . 
Er gruppledare får era valsedlar . 
Ni markerar era valsedlar som er ledare och visar dem för observatören . 
Är det så svårt ? 
- Okej , då ska vi se . - Hej . Mobiliseras verkligen regeringsarbetare ? 
Ja , men det slutar inte där . 
Vi fick tips om att de övade på att rösta . 
- Övade ? - Ja . 
De övade på att rösta på president Rhee . 
- Vet du var ? 
- Ja , ska jag åka dit ? 
Ja , åk dit och ta reda på mer . 
Ja , herrn . 
Nästa . 
En uppföljning av Kang Seongmin och Sineuialliansen . 
Kopplingar mellan Sineuialliansen och Kang Seongmin 
Vi släpper det . 
Misstankarna kvarstår ... 
Låt det vara . 
Nästa . Berätta vad du fick reda på . 
Ja , herrn . 
Vad är det ? 
Journalister som skrev om Sineuialliansen blev utpressade . 
Chefen tänker bara på ditt bästa . 
Enligt polisrapporten sköts Yoon Palbong först . 
Även andra skottet var riktat mot honom . 
Vad betyder det ? 
Jag vet inte . 
Ska vi bara låta det vara ... med alla obesvarade frågor ? 
Jag ska prata med inspektören som hanterade Sineuialliansen . 
Kapitalförsvarskommandot 
Lägg dem här . 
Vad är det här ? 
Det är gåvor , herrn . 
Gåvor ? 
Jag beställde dessa åt dig från en affärsman som importerade varor till logistikkommandot . 
Har ni hittat några Sineuialliansmedlemmar ? 
Varför svarar ingen ? 
Välkomna , polischefer . Koreas framtid hänger på det kommande valet . 
Låt oss samarbeta för att skydda vårt land . 
Låt oss skydda Korea ! 
- Skydda det ! - Skydda det ! 
- Låt oss vinna ! - Låt oss vinna ! - Låt oss vinna ! - Låt oss vinna ! - Låt oss vinna ! - Låt oss vinna ! 
Arméns Counter Intelligence Corps 
Hong Youngki kan märka vem som helst som kommunist . 
Hur ? 
Han kokar ihop bevis och burar in dem . 
- Fånga kapten Kim först ! 
- Vad händer ? 
Han sparkade en tredjedel av generalerna . 
Släpp ! 
Vägen till samexistens Inte ens en general kan göra mycket under hans uppsikt . 
- Ta honom ! 
- Få ut honom nu ! 
- Stanna inomhus , barn ! 
Era jävlar ! 
- Kom hit ! 
- Vart för ni mig ? 
Vad händer ? 
- Släpp ! - Rör på er ! 
- Pak Wonil . 
- Ja , herrn . 
Känner du till Arbetarpartiets 29:e direktiv ? 
Nej . 
Arbetarpartiets 29:e direktiv . " Infiltrera armén - och vinn över högt uppsatta . " - Nej . 
Jag har aldrig hört det . 
Ta en cigg . 
Det friskar upp minnet . 
Hej då ! 
Vilka är ni ? 
Varför står ni i vägen ? 
Vi är från åklagarmyndigheten . 
Åklagarmyndigheten ? 
Och ni har fräckheten att stå i vägen för en ledamot ? 
Ta honom . 
- Håll fast honom . 
- Släpp ! Jag tar Pak Jiwook med Han Soo som lockbete . 
Och sen ? 
Sen tar jag Choi Hanrim med Pak Jiwook . 
Hong Youngki har planterat bevis . 
General Min Soochul kommer att gripas för spionage . 
Vi hittade den i din vas . Förklara . 
Jag har redan mutat kapitalförsvaret . 
Jang Doosik blir befälhavare för kapitalförsvarsenheten och Jeong Hanmin vice befälhavare . 
Vice befälhavare Jeong Hanmin till er tjänst . 
Då hamnar Choi Hanrim i Jang Doosiks och Jeong Hanmins våld . 
Tack , befälhavare Jang . 
Hej . 
Här . 
Adresserna är fem år gamla , så de kan ha flyttat . 
Tack , herrn . 
Varför granska alliansen ? 
Cha Taemin har inte fångats . 
Vi försöker inte ens . 
Saknar Kang Seongmin koppling till alliansen ? 
Ledamot Pak Jiwook tog nyligen deras adresser . 
Han samlade tidigare underhuggare från Folkets fredsbyrå . 
Ledamot Pak Jiwook ? 
Sluta be mig om tjänster . 
Det är hektiskt även för polisen som mobiliseras . 
Mobiliseras polisen ? 
Har du officiella dokument på det ? 
Nu räcker det . 
Vad är det med dig ? 
Lista över Sineaualliansens medlemmar 
Ledamot Pak Jiwook rekryterade före detta poliser . 
Att skugga dem kan leda dig till Cha Taemin . 
Varför skulle ledamot Pak göra det ? 
Det känns som om Kang Seongmin är inblandad . 
Val påverkade av regeringsmanipulation , mutor och olagliga aktiviteter ... 
Varje tecken på korrupt demokrati uppenbaras framför våra ögon . 
Demokrati 
Med maskopi , konspiration och skenhelighet ... 
Tack . 
... verkar valet bli än mer förvirrat . 
Oavsett vem som vinner , kommer kaos att uppstå . 
Eftersom politiker är upptagna med sina egna maktkamper , får vi se om detta politiska kaos ... 
Tack . 
... blir Koreas växtvärk eller dödsdom . 
Från och med nu är Sineuialliansen återinsatt . 
Vi kämpar mot auktoritet , makt och orättvisa . 
Intellektuella har sålt ut sitt samvete , politiker sin ideologi och folket sitt hopp i vår tid . 
Medvetna medborgare måste resa sig . 
Det är svårt att återta det som har tagits ifrån oss . 
Ingen kan kämpa för oss . 
Demokrati betyder att suveränitet tillhör folket . 
Vem ska skydda det som är vårt om inte vi gör anspråk ? 
Sineuialliansen är beväpnad och kämpar mot orättvisor . 
Sineuialliansen står upp mot den makt som förtrycker vårt folk . 
Vi motsätter oss allt och alla som monopoliserar makt och är beredda att använda våld och vapen . 
Alla som förespråkar förtryck ska straffas i Sineuialliansens namn . 
Okej , uppfattat . 
Farbror Samsik . 
Oroa dig inte . Det lugnar ner sig . 
- Vi är studenter ! - Kan du få studenterna släppta ? 
- Givetvis . 
Och kaptenerna Kim Inho och Pak Wonil ? 
De hålls på CIC . 
De erkänner i morgon bitti . 
Jag vill erkänna nåt . 
Vad är det ? 
Jag låg med Rachael . 
Det förklarar ditt goda humör . 
Jag slutar om du ber mig . 
Tänk på Rachael ... som en blåsfisk . 
När giftet är borta kan den bli en utsökt rätt . Men om giftet finns kvar kan det vara dödligt . 
Statskuppen var hennes idé . 
Jag vet . 
Kan vi fullfölja vår plan ? Ja . 
Vi behöver bara följa planen . 
Tänk om det går snett ? 
Livet går ofta snett , men man blir aldrig fri från sina planer . 
Vem kan vi skylla på ? 
Det är bara så livet är . 
