Vi hittar Chimera och dödar Chimera . Enkelt . 
Så vi ska till kusten ? 
För femtioelfte gången , det var där varelsen var . 
Den har såklart flyttat till klipporna nu . 
Vet du vad ? Jag är så trött på att du ifrågasätter mig . 
Om du inte var så kortsynt ... Ursäkta , " kortsynt " ? 
Driver du med min längd ? 
Nej , med din tjocka skalle . 
Det räcker nu . 
Vi delar på oss och letar efter spår . 
Ni kan väl gå ihop ? Ni har ett så unikt förhållande . 
Underbart . Barnvakt igen . 
Ja , ja . Håll jämna steg , spända jävel . 
Som jag sa , vid kusten . 
Du menar klipporna nära kusten . 
- Kima , vänta ! 
- Jag klarar det . 
Det gör du inte . 
Allura ! 
Kima ! Ducka ! 
Försöker du ta livet av dig ? 
Ur vägen , sa jag ! 
Jag sa ju att jag klarar det . 
Kima ... 
Var är du ? 
Skit . 
Nåt ? 
Vorugal är kvar där nere . Jag känner det . Vad väntar vi på då ? 
Vi kan inte ge oss på en drake utan en plan . 
Planen är att jag hittar Kima och sliter det jävla monstret i bitar . 
Strategin har några fördelar , men vi är för få för ett drakanfall . 
Och vi har ont om tid . 
Om en timme måste vi öppna porten åt våra vänner . 
Varför plötsligt så försiktiga ? 
Skulle du vänta om Vex ' ahlia var i fara ? 
Skulle du avvakta om Percivals liv hängde på en skör tråd ? 
Det är fullständigt ... 
Percy och jag är inte ... Ni är inte vad ? 
Vi är inte ihop . 
Ni hade kunnat lura mig . 
Men du har en poäng . 
Vi har alltid gett oss in i fara för varandra . 
Det vore hyckleri att inte göra det nu . 
Tack . 
Det var det jag menade . 
Att vara ihop skapar alla möjliga komplikationer . 
Men vi är väl inte ihop ? 
Va ? 
Nej . 
Då är det inte komplicerat . 
Jag undrar hur det går för de andra . 
Säkert bättre än för oss . 
Varför är det så djävulskt långt till porten ? 
Tror du att du kan ta oss , dingelsnorre ? 
Du kanske inte ska håna mördarmannen . 
Jag vet att du är där . 
Det är bara en tidsfråga . 
Fortsätt gömma dig , råtta . 
Jag hittar dig . 
Märkligt . 
Isen där nere ser tunn ut . 
Vi kan dra nytta av det . 
Strunta i isen . Ser du Kima ? 
Fotspår ? Nånting ? Inte härifrån . 
Då går vi närmare . 
Ha tålamod . 
Vi ser inte draken . 
Det är Kima . Hon har inget tålamod . 
Utan mig försätter hon sig i större fara . 
Vi kanske ska följa Allura . 
Jag har aldrig sett henne så impulsiv . 
Desto viktigare för oss att behålla lugnet . 
För vi är alltid så förnuftiga . 
Har kylan börjat påverka dig ? 
Fan ta det här . 
Spring , lilla hare . 
Som du vill . 
Där är hon ! 
Jag har dig nu . 
Kima ! Här borta ! 
Allie ? 
Fan . 
Håll ut ! 
Perfekt . 
Vänta . Förnuftiga , minns du ? 
- Tog en . 
- Ner ! 
Vad fan , Allie ? Gå undan . Jag klarar det ! 
Bevisen talar emot dig . 
Nej ! 
Ja ! 
Kom igen , slå tillbaka . 
Håll det intressant . 
Förnuft fångat . 
Snyggt skott . 
Jag hittar Kima . 
Möt mig vid portalen ! 
Vill du ha en utmaning ? 
Fan ta mitt liv . 
Vilken härlig , bottenlös grop du har hittat , älskling . 
Ganska rymlig . 
Tack för att du fångade mig . 
Kan du få ut mig ? 
Ledsen . 
Fenthras har en egen vilja ibland . 
Ditt vapen är jävligt högljutt ! 
Ledsen , alla kan inte skjuta magi ur fingrarna ! 
Jösses . 
Percy ? 
Han verkar ha övergett dig . 
Har jag ? 
Det är långt ifrån över . 
Skit . 
Dags att improvisera . 
- Förlåt , jag lyssnade inte ... 
- Glöm det . Vi letar upp våra kvinnor . 
Var fan är porten ? 
Jag vet inte ! Klipporna ser likadana ut ! 
Den borde vara rakt fram . Den är bara stängd . 
Nåt måste ha hänt de andra . 
Keyleth , kan du öppna portalen härifrån ? 
Jaså ? Låter svårt . Försök ändå ! 
Där är den ! 
Jag kan börja . Men de måste aktivera den på andra sidan . 
Tror du att han ger oss fem minuter om vi frågar snällt ? 
Antagligen inte ! 
- Allie . - Kima ! 
Vad fan tänkte du ? 
Jag sa åt dig att låta bli . 
Så du kunde kasta dig in i Vorugals käft ? 
Nån måste rädda dig från dig själv . 
Jaså ? Det igen ? 
Varför kan du inte lita på mig ? 
Jag ... Jag kan inte ... Du är oberäknelig och det skrämmer mig . 
Förlåt . 
Jag gör inte det här för att jag har en dödslängtan . 
Det är bara ... mitt sätt skydda dig . 
- Tjejer ? 
- Porten . 
- Ja , förestående undergång . - Ja . 
Inte min styrka , men jag försöker . 
Nej ! 
Han har hittat oss . 
Vi behöver mer tid . 
Vi håller honom ute . 
Eller inte . 
Stoppa honom så länge ni kan ! 
- Vax , är du galen ? 
- Det verkar så . 
Hörni , Vax är i trubbel ! 
- Ja . - Vi hämtar honom . 
- Åh , gud . 
- Scanlan , nu ! 
Toppen . Nu är jag också galen ! 
Grog . 
- Kiki ! Nåt ? 
- Den rör sig inte ! 
Eld . 
Jag kanske kan absorbera den ! 
Pike ? Pike ! Gå därifrån ! 
Skölden ... Jag tror att det fungerar ! 
Jäklar ! 
- Fan . Ditt huvud ! 
- Vad är det med det ? 
Vad fan ? 
Hörni , titta ! Portalen ! 
Skit , jag vill inte dö skallig ! 
Rör på er ! 
Kom igen ! 
Ja ! Det är dem . 
- Hjälp , hjälp ! 
- Stor , stor kille jagar oss ! 
Fan ! 
Vad är det för grej ? 
Tror du att de kommer att slåss eller knulla ? 
En demon mot en drake ? 
Jäkligt grym plan . 
Det är det vi är kända för . 
- Pike , ditt hår är ... 
- Käften , de Rolo . Jag har en dålig dag . 
Flyg ! 
Herrejävlar . 
Alla till mig nu ! 
Vänta , vänta ! 
Okej , kör ! 
Den här uppvisningen är fantastisk ! 
Ja , för fan ! 
Okej , fem guld på eldkillen . 
En en-två-kombo . 
Ta honom . 
Slår på stort ! 
Såg du det ? 
Vi kanske ska kolla därifrån . 
Ja , lite avstånd låter bra . 
Ur vägen ! 
Du förlorar . 
Är det över ? 
Han kanske är för trött för att slåss . 
Varför måste ni utmana ödet ? 
Ja , du har rätt . 
Förlåt . 
Vad ska vi göra ? Fly ? Attackera ? 
Jag har en idé . 
Vänta här . 
Va ? 
Hallå , den är min ! 
Vart fan ska hon ? 
Oroa dig inte . 
Det är lady Kima av Vord . 
Bestmördare , överlevare av Emberhold , och kvinnan jag älskar . 
Hon klarar det . 
Ja , kom . 
Okej . Lite hjälp nu . 
Du hörde henne . 
Vi har dig , Kima . 
Sätt igång ! 
Han ger sig av ! 
Titta vad jag fångade . 
Jag tänker inte hållas fast ! 
Hur kan den fortfarande leva ? 
Jag vet inte . Det är en drake . 
- Kan du förtrolla ett rörligt mål ? 
Kima ! Är du fortfarande med mig ? 
Dö , byte ! 
Tack , älskling . 
- Redo ? 
- Nej , men gör det ändå . 
Var försiktig med vad du jagar . 
Än en gång ger du dig in oavsett faran . 
Det är ... okej , va ? 
Det var det jag föll för . 
Kom hit , din spända jävel . 
Jag vet . Vi är inte ihop . 
Men vi behöver inte vara åtskilda . 
Drakfjäll . 
Vorugal . 
Ännu ett misslyckande . 
Värdelösa , allihop . 
Alla är emot mig , men det kvittar . 
Min avkomma kläcks . 
De behöver bara sitt första byte . 
Är det så ? 
Vem är det ? 
Jag har det perfekta stället i åtanke . 
Hår . 
Vilken lättnad . 
- Inget illa menat , kompis . 
- Ingen fara . 
Inte många kan bära upp den stilen . Om du förstår ? 
Det blir mörkt snart . 
Allura , kan du " bamfa " ut oss härifrån ? 
Jag måste tyvärr vila innan jag kan " bamfa " nåt . 
Vi kan ta in på slott Shorthalt . 
Var ? Ni vet , mitt vattensängshem ? Det heta stället . 
Shortkåken . Ni vet , min nattklubb . 
Vi är för trötta för skämt , Scanlan . 
Tro mig , ni skulle skratta om jag skämtade . 
Jag kan inte göra det utan en dörr . 
Menar du så här ? 
Grog , du är fantastisk . 
Okej , jag stoppar in min magiska nyckel och ... 
Scanlan , vad fan är det ? 
