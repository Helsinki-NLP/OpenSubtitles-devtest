- De har dödat domaren ! - Kom igen ! 
Låt dem inte komma undan ! 
Vad hände ? 
Jag är inte tränad för det här . Det var vad som hände . - Jag trodde att jag skulle stupa först . - Ja . Samma här . 
- Det kommer fler . 
- Vi kommer inte förbi dem . Vi måste . Det är enda vägen hem . 
Kanske inte . 
Bärarna ? Har du med dem att göra än ? 
Vi måste ta oss ner två nivåer till . 
Försök att hänga med . 
Det är så uppenbart att det var du . 
Varför då ? 
Han vet inte namnen på mina lyssnare , men han ser kännetecknen . 
Han spårade kampanjen för att avsätta Meadows tillbaka till mig . 
Mamma . Mamma . - Ett ögonblick , vännen . - Det är en man i köket . 
Kan jag hjälpa dig ? 
Jag minns inte när jag lagade mitt eget kaffe senast . 
Jag talar sällan om borgmästare Jahns , men hon lagade jämt sitt eget kaffe . 
Hon sa att vardagssysslor som vanligt folk i Silon ägnar sig åt hjälpte henne att känna en koppling till dem i brist på annat . 
Ni förstår , det här jobbet kräver att jag har ett annat perspektiv än nån annan . 
Låt mig göra det . Maskinen är knepig . 
Jag är känd för att vara bra på maskiner . 
Du jobbade med Rob förut , va ? 
Jag jobbade för honom , som han gärna påminner mig om . 
Diskuterar han jobbet med dig ? 
Robert vet att jag inte är så intresserad av det jobbet mer . 
Jag har mitt jobb hos IT och min son . 
Pakten säger : " Mödrar är ett kärl för att föra våra barn till världen , liksom Silon är ett kärl för folket . " 
I vår familj tar vi allvarligt på det . 
Er familj läser Pakten tillsammans , berättade du visst ? 
Varje kväll . 
Kan du hämta ert ex av Pakten åt mig ? 
Visst . 
Du svek mitt förtroende , Rob . 
Du tvingade mig att göra nåt jag inte ville göra . 
Du är inte längre säkerhetschef för Rättsavdelningen . Du kommer inte att bli min skugga . Men du är för värdefull att avvara helt . Så du får ta Marys jobb . Du ska bli domare . 
Lägg din hand på Pakten och upprepa efter mig . 
Jag , Robert Sims , svär högtidligt ... BASERAD PÅ BOKSERIEN SILO AV HUGH HOWEY 
Jag ska ta en titt . 
- Är Calvin här ? - Vem är det som frågar ? 
Calvin . Det var ett tag sen . 
Jag slutar alltid att se bärare efter en viss ålder . Knäna . 
Ska en kvinna i din ställning börja med en förolämpning ? 
Var glad om nån del av dig klarar sig tillbaka ner . 
Det är därför vi är här . 
Vi behöver en plats att vila på , och jag behöver transport hem för mig och mina vänner . Det är inte gratis . 
Möjligen har jag en låda av bourbon från tiden före . 
Det kostar mer än gammal sprit . 
Har du nåt som tillhörde Juliette Nichols ? 
Hej . Vad gör du ? 
Tja , jag fick ingen brandmanshjälm , och jag vill inte gå ner i vattnet igen . Så jag prövar om min gamla funkar . 
Du , jag tänkte fråga en sak . Er generator är hundra nivåer under vattnet . Så hur kan lysena vara på ? 
IT har sin egen kraftkälla . 
Den kommer utifrån . 
Utifrån var ? Där uppe , typ ... Vet du varför generatorn slutade fungera ? 
Jo , några soldater från Rättsavdelningen fick den ljusa idén att spränga länspumpen på 144:e för att spola ut Mekaniska . Men de hann inte laga den innan vattnet kortslöt generatorn . Så vattnet fortsätter ... Jag förstår . Finns det ... Finns det ett sätt att få vattnet att sluta stiga , tror du ? 
Den närmaste länspumpen är på nivå 30 . Under vatten . Men man kan dra elkraft till den . Kanske hindra att vattnet stiger mer . - Ja . - Vänta , du ... 
Du kan stoppa det . Jag ? Nej . - Hinner inte . Jag måste göra det här . - Jag har inte tid . - Tiden rinner ut för mig . - Inte alls . - Du har månader , år att tänka ut ... - Tio månader . - Jag har tio månader . - Tio månader ? Jag har dagar . Men det kan du inte veta säkert . 
Så varför ska jag ta risken ? 
Om tio månader rinner vattnet in i IT . 
- Om 13 är det helt under vatten . - Nej . Sluta ! 
Det här är vad jag måste göra . Och den där funkar inte . Okej ? 
- Den går inte att koppla in . - Vart ska du gå ? Jag måste ta mig till dräktrummet för att hitta en hjälm som funkar . 
Hallå , vänta ! 
Var är de ? 
De lämnade trappan på nivå 70 . Kameror slocknade och vi vet inte var de är , men jag skickade soldater . 
De är förklädda till civila och uppviglar mobbar från 60:e ner till 130:e . 
- Satte du pris på ledarnas huvuden ? 
- 1 000 krediter var . Be Rättsavdelningen sätta upp barrikad på 130:e , ifall de kommer undan . 
De kommer inte förbi mitt folk . 
Gör mig till viljes , mr Amundsen . Jag oroar mig . Det är mitt jobb . 
Och eftersom vi har bråttom ska jag ignorera att du sa " mitt folk " . 
Låt mig vara tydlig . Rättsavdelningens soldater är på intet sätt " dina " . 
Vi fick just meddelande . De befinner sig på 70:e . 
Hur vet jag att det är hennes ? 
Det vet du inte . Men jag vet . För jag gav det till henne för 20 år sen . 
Och jag lagade gångjärnet när hon försökte bända loss fastfrysta bultar , vilket jag avrådde henne från . 
Jag tar den . 
Plus de 24 kylspolarna du utlovade för din vistelse här . 
Släng med den fina spriten , så är vi överens . 
- Vad är din plan ? - Sädesbingar . 
Alla vet att kvarnen på nivå 59 fallerar varannan vecka . 
Ingen kommer att bevaka säd på väg ner till de lägre nivåerna . 
- Fan heller . - Jag sa inte att det blir bekvämt . 
Jag pratar inte om bekvämlighet . Men vi har en fjärde person . Rätt stor . Han får aldrig rum . 
Det är enda sättet . 
Nedstigningsriggen , då ? 
- Vet inte vad du menar . - Jodå . Inte jag . 
- Ett system med eldriven vinsch . 
- Det strider mot Pakten . Och du fixade den i enlighet med Pakten ? 
Vi tog den ur cirkulation , bara . 
Bärarna har ensamrätt att forsla gods i Silon . 
Om folk ser det där , börjar de få andra idéer . 
Vi måste iväg ! Soldaterna kommer . Fort ! - Du meddelade Rättsavdelningen ! - Jag tänkte hjälpa er . Men en belöning är utfäst . Den är för hög att ignorera , även för gamla vänner . 
- McLain ! - Den jäveln ! 
Enligt Doc Phelan har inte Kennedy varit hos honom . 
Kennedy kanske känner hans rykte . 
De bästa får jobb på Toppnivån , vi får ta de som blir över . 
Frånsett mig , förstås . 
Vad är det ? 
Ett meddelande från Rättsavdelningens nya chef . 
Rick Amundsen . 
Sims , då ? 
Han är insatt som domare . 
Var är Meadows ? 
Död . 
Mördad . 
Va ? 
Av chefen för Mekaniska och hans kollega . 
Knox och Shirley ? 
Det där liknade inte Jules multiverktyg . 
Nej , det var mitt . Jag vet inte var hennes är . 
Försiktigt . Jag har dig . - Okej . - Gick det bra ? Bäst att vi delar på oss , så vi inte saktar ner er . 
Belöningen gäller oss två . 
Alla löper risk att bli dödade . 
Bli inte gråtmilda nu . Stick . Gå . 
- Du följer inte med . 
- Va ? Du kanske inte förutsåg det här scenariot när du stängde in dig i din verkstad för 25 år sen . Men nu vet ingen över nivå 125 vem du är . 
Det är din smala lycka . Jag , däremot , är chef för Förrådet . 
- Carla , jag vägrar ... - Martha . 
De behöver dig där nere . Nu mer än nånsin , troligen . 
Gå . 
Bara ett vanligt skrubbsår . 
Rengör det med tvål , så läker det fint . 
Får jag se . Okej . Det är inte så farligt . Tryck på såret , bara . 
Jag är strax tillbaka . Nejlikolja hjälper mot värken , och det väldoftande hjälper dig att sova . 
Tack . Det doftar gott . Det knäppte till i axeln . Jag behöver läkare . LÄKARSTATION Bra idé . Han är där borta . 
Fan , vad ont det gjorde . 
Rör på axeln . 
Ja . Glöm inte nejlikoljan . - Tack . - Ja . 
Imponerande teknik för nån som bär på en bebis . 
Tack . Min mor var örtkännare . Och pappa var ett fyllo som förlorade många slagsmål . Dr Pete Nichols . 
Angenämt . 
Kathleen Billings . Som i sheriff Billings ? 
Jag förstår varför du är här och vårdar skadade . Det skingrar tankarna . 
Jag kan inte sitta hemma . Jag blir nervös . 
Paul skickades till Mekaniska . Det var nån incident där nere . 
- Jag hörde om det . Nån brand eller ... - Dr Nichols . 
Ja ? Följ med oss , tack . 
Nu . 
Vad är hans plan ? 
Låta Silon ta hand om mördarna . 
Om han lyckas blir det som en nystart för honom . Som om det där med Juliette Nichols aldrig hänt . 
Du har gjort såna uppdrag . Civilklädda soldater . 
Stor belöning för rymlingarna . Låt mobben jaga dem . Kanske ta lagen i egna händer . 
En sån känslig operation kräver erfarenhet , Rob . 
Amundsen är bra . Han har haft bästa tänkbara lärare men är inte bäst . 
Tänk om han inte klarar det ? 
Gör det bästa av jobbet , Robert . 
Dr Nichols . Tack för att du kom . 
Om du tror att jag vet nåt om de där från Mekaniska , har du fel . 
Nej då . Nej . Nej , det har inget med det att göra . 
Jag tänkte att du ville ha några av din dotters saker . 
Vanligtvis skulle dessa saker återanvändas , men dessa omständigheter är långt ifrån normala . 
Om dessa saker återanvänds , är jag rädd att de skulle vördas , åtrås , skapa avund , oenighet och slutligen våld . 
Det vore inte enda sättet på vilket din dotters minne har förvrängts för att passa andras agendor . 
Jag hörde att du vårdade folk som skadats i upploppet efter mordet på domare Meadows . 
Den tjänstvilligheten ger mig hopp om att du kan vara en viktigare del av denna rörelse . Rörelsen för att återställa ordningen i Silon , och tron på Pakten . 
Och om jag säger nej ? 
Varför skulle du säga nej ? 
Jag vill bara ha klarhet . 
Om jag inte hjälper er , vad händer då ? 
Jag har inget kvar att mista , eller hur ? 
Silon har tagit min son , min fru och nu min dotter . 
Jag vårdade inte skadade av plikttrogenhet mot Silon . Jag försökte bibehålla min yrkesmässiga integritet . Jag försökte praktisera sjukvård utan lögner , utan skada . 
Och de där fejkade borttagningarna av födelsekontroller ... Jag ser de där unga paren . Deras ansikten lysande av hopp . Hopp som jag vet är ogrundat . 
Mitt yrke är bluffmakeri . 
Silon tog det också från mig . 
Hursomhelst är min dotter död . Du kan inte styra över vad hon betyder för folk . Eller vad hon betyder för mig . 
Så , Solo ... - Ja . - ... är det ditt riktiga namn ? 
- Co ... Cole Myers heter jag . 
- Cole . Jag gick på en tillställning och de frågade : " Vem är du med ? " Jag sa : " Jag är solo " , och Russells grabb var där och hörde mig säga det , och trodde att det var mitt namn , så jag fick heta det . 
Men alltså , vad betyder ett namn ? 
Okej . Det är från din pjäs . Romeo och Julia innan de dör . 
Innan vilka dör ? 
Romeo och Julia . 
- De dör inte . Nej . - Jo , det gör de . I vår pjäs dör de . 
- Helvete . - Är du okej ? - Jadå . - Är du hungr ... Jag vet inte , jag är bara ... trött . Jag är okej . Är du hungrig ? 
- Vet inte . Ja , kanske . 
- Ja ! - Okej , men ... - Jag ska gå och hämta mat . 
Helvete . 
RÄTTSAVDELNINGEN Ni får kopior av de här rapporterna . 
Om de har små flaggor , följer rekommendationer från borgmästarämbetet . 
När ni har nått ert beslut , - skriver ... - Jag har varit här i många år nu . 
Visst , domaren . 
Vi har ännu inte kunnat fabricera din signaturstämpel . Så om du kan underteckna tills vidare ... Domare Sims ? 
Bra jobbat . 
De andra ? 
De två med belöningar på huvudet är i trapporna . 
Jag har civilklädda soldater några nivåer längre ner . Och vi uppviglar mobben . 
Säg till när ni har gripit dem . 
Ska bli . 
Tack , du kan gå . 
Mr Kyle . Hur är det nere i gruvorna ? 
Det har bara gått en dag . 
Du lever än i alla fall . Det är bra . 
Vet du hur länge folk överlever i genomsnitt där nere i gruvorna ? 
Nej , sir . 
Fem år . 
Så när domare Meadows halverade din dom , var det på sin höjd en symbolisk gest . 
Det är inte troligt att du överlever din tid där . 
Vet du varför ? För att det är farligt ? Gruvras , kvävning , krosskador , mista armar och ben , sprängningar som gått fel . 
Det är hård regim . 
Jag ska erbjuda dig lite lätt regim , Lukas . 
Jag har ett projekt där din hjärna behövs . 
Dagen då domare Meadows mördades berättade hon att du kunde ta små spridda bitar information om ljusen på natthimlen och skapa en modell som , oss emellan , var ganska exakt . 
Stämmer det ? 
Jag har en annan sak som består av fragment , och som jag vill att du rekonstruerar . 
Känner du igen den ? 
Det är hårddisken som Juliette Nichols visade dig . 
Du kan säga som det är . 
Du kommer inte att straffas för det . 
Ja , jag känner igen den . 
Jag krossade den , för den är en förbjuden relik som troligen innehåller farlig information . 
Men jag har inte längre råd med ovetskapens lyx . 
Du måste ta reda på vad som finns på den . 
Du kan jobba härifrån . 
Har du några frågor ? Kom igen nu . 
Du vet säkert att det finns minst tre personer där ute i IT:s pool som klarar det här bättre än du . Men jag vet att du kommer att jobba hårdare än nån jag kan hitta där ute för , tja du vill leva längre än fem år . 
Domaren , är allt som det ska ? 
Säg det du . 
Knappen fungerar inte . 
Vi har allt i ordning här , Ers nåd . Ers nåd ? Domaren ? 
Säg Rob som du har gjort de gångna tio åren . 
Jag försöker räkna ut det här , precis som du . 
Jag var nyss i mitt kontor . Mitt nya kontor . 
Jag satt bakom samma skrivbord som kvinnan jag jobbat åt i 15 år . Det vore en bra idé att se hur det går med sökandet efter dem som mördade henne . 
Jag ska ordna att du får alla relevanta detaljer imorgon bitti . 
De misstänkta är kvar i trapporna . 
Vi använder planen du beslutade om . 
Fortare . 
Värst vad du har bråttom . 
Hej , min man och jag är på väg ner för att träffa några vänner . 
Det verkar oklokt . Farliga mördare på fri fot . 
Och vad gör ni ute ? 
- Vi är bekymrade medborgare . 
- Och vem är du ? Få se legitimation . 
Kräver Pakten att medborgare identifierar sig för andra medborgare , vare sig bekymrade eller ... 
- Nej . - Nej , den ... Han är beväpnad ! 
Sluta ! 
Sluta , sa jag ! 
Några känner visst igen mig . Och jag känner igen några av er . 
Ni vet vem min man är . Men ni kanske inte vet om hans nya position . 
Domare Sims vill att de här rymlingarna grips . 
Vill ni döda dem här och nu ? Det vill jag också . Men rättvisa för domare Meadows är inte bara vår sak , utan en sak för hela Silon . 
Och alla kommer att se på när de här två går ut för att putsa . 
Följ med mig , annars kommer ni att bli lynchade . 
Fan också . 
Här är ni säkra så länge . 
Tar du oss inte till Rättsavdelningen ? 
Kamerorna funkar än i trapporna , men här är de trasiga . 
När de ser mig gå upp ensam skickar de fler soldater efter er . Kanske många . Så vänta ett tag innan ni går . 
Det finns en barrikad på 130:e . 
Jag vet inte hur ni ska ta er igenom , men det är ert problem . 
Varför hjälper du oss ? 
Camille . 
God morgon , Asa . 
Du går till jobbet tidigt idag . Och du blir hos din exfru ikväll , på 83:e . 
- Jag slutade nyss nattskiftet . 
- Då kommer din chef att tänka att du är den flitigaste rörmokaren i Silon . 
Ge mig nycklarna . 
Vad i helvete , Camille ? 
När du får höra om en belöning för dem som mördade Meadows ignorerar du den , så fortsätter jag ignorera dig . 
Förstår du ? 
Låt mig åtminstone ta på mig byxorna . 
Varför tog du inte på dig dem först ? 
PAKTEN MELLAN GRUNDARNA OCH SILONS MEDBORGARE Är de infångade ? 
En rätt stor konflikt , va ? 
Vadå ? 
Att vara vicesheriff när mina vänner jagas som mördare av halva Silon . 
Nästan lika stor som att lova att genomdriva Pakten och samtidigt ha en sjukdom som uttryckligen fördöms av Pakten . 
Vet de ? 
Sims vet . 
Som chef för Rättsavdelningen lät han det passera . Som domare ... Jag kanske vet var Patrick Kennedy är . 
Försök att inte äta upp allt i kylen . 
Jag är bara en hårt arbetande kille vars huvudjobb är att hålla Silon igång . 
- Det beror på vad som finns där . 
Jag bara skojar . 
Hur tror hon att du ska komma in utan nyckel ? 
Det tror hon inte . Om hon vill att jag ska ha den , får hon den till mig på nåt sätt . 
Ett gott råd , stanna så länge ni behöver . Men stick innan hon är tillbaka . 
Jag hjälper henne inte av artighet . 
Jag gick med på det för att jag är rädd för henne . 
Det borde ni också vara . 
Han bor för fan i en garderob . 
Tror varje avdelning att det är just de som håller Silon igång , tror du ? 
Förmodligen . 
Jag har sagt samma sak för att samla alla i Mekaniska . 
Det fungerade för att det är sant . 
Även om resten i Silon tror nåt annat . 
Du är en bra ledare , Knox . 
Mekaniska hade gått åt skogen för länge sen om det inte var för dig . 
Jag hade fel om taktiken . 
Jag ville be vänligt ... Nu måste vi dö för det . 
Vi hade aldrig en chans från början . 
Men om vi hade gjort på mitt sätt hade vi redan varit döda . 
Tror du att Knox och Shirley dödade domare Meadows ? 
Uppriktigt ? Sen Jules gick ut har allt gått överstyr . 
Shirley och en mobb angrep min station . Nu har Knox lierat sig med henne . De saknar respekt för ordningen i Silon . 
Tror jag att de dödade Meadows ? Inte en chans i helvetet . 
Vänta lite . 
Frances . Vänta lite . Vart ska du gå med den där maten ? 
Hem ? 
Det är efter midnatt . Ditt skift började kl 06 : 00 . Så istället för att sova stannar du uppe och äter samma mat som du har serverat i 18 timmar ? 
Såvida det inte är förbjudet , Hank , så är det vad jag gör . 
Vi kan din historia , Frances . 
Doris Kennedy var din faster och du sålde piller som hon stal . 
Har du bevis ? 
För det hade du inte för fem år sen . Lugn , Franny . Vi är inte här för det utan för att vi tänker att din farbror Patrick inte kan leva länge till bara på varma måltider . 
Så låt oss ta med maten , vetja . 
Hur var din första dag , domare Sims ? 
Jag skrev på där de sa . 
Jag gick till Bevakarnas rum för att få fakta om mördarjakten . 
Amundsen släppte inte in mig . 
Men han sa att tre av de misstänkta ännu är på fri fot . 
Om du var chef hade de varit gripna för länge sen . 
Ursäkta mig . 
Jag bor i 132 . 
Inte ikväll . 
Jag jobbar hos polisen . Vi blev inte informerade om det här . 
Det här rör inte polisen . 
Om Rättsavdelningen tror att de kan utestänga medborgare ... Vänd och gå tillbaka samma väg . 
Skojar du ? 
Ni har ingen rätt att konfiskera lägenheten för en polisanställd . 
Jag måste ... Så fort vi är i trappan ser de oss . Och så fort vi stänger dörren är vi utelåsta . 
Vi måste gå hem nån gång . Vi tar trapporna och springer som fan . 
Okej . Men inte nedåt . - Uppåt . 
- Va ? 
Lita på mig . 
JAY , SUNIL LÄGENHET 101 , NIVÅ 16 PENN , MARJORIE LÄGENHET 57 , NIVÅ 23 SAMUEL , TRINA NIVÅ 17 , KORTNAMN : TINY De fastnade i folkmassan . En f.d. soldat gömde dem på 73:e . Vi kollade varje lägenhet . Inget resultat än , - men jag har stängt sopnedkastet . - Vänta lite . 
Varför gömde en f.d. soldat dem ? 
Hon var rädd att de skulle lynchas . Vem var hon ? 
Camille Sims . 
Hitta de där jävlarna från Mekaniska . 
- Hur långt upp ska vi ? 
- Håll tempot bara . 
Jag lyckades bara rädda några saker . 
Jag fann några fragment som överlappar filer i vår databas . 
Här är vår karta över Silon , och jag har använt denna fil för att fylla i lite saknad data från ett av fragmenten , som också är en karta . 
Den skiljer sig från vår karta över Silon på några ställen . 
Det finns linjer som kommer från utanför Silons väggar . Det finns nåt på IT-nivån och nåt på Rättsavdelningen . 
Nån aning om vad det är ? Nej . Det finns nåt mer . - Där , på själva botten av Silon ... - Vad är det ? 
- En tunnel . 
- Vart leder den ? 
Jag har ingen aning . 
Nåja , fortsätt jobba . 
Du har tjänat ytterligare 24 timmar utanför gruvan , mr Kyle . 
Sir , det fanns också en mapp som jag hittade . 
Jag kunde återskapa den oförstörd , och de flesta filerna var bara PM från avdelningarna , men en var annorlunda . 
Det var en skanning av ett handskrivet brev till nåns hustru . 
Vem ? 
Salvador Quinn . 
Vad stod det i brevet ? 
Det är ett kärleksbrev , men sen blir det lite konstigt . 
- Det övergår i , typ ... - I kod . 
Ja , just det . 
FARA ! ATT FORTSÄTTA LÄNGRE ÄR ETT STRAFFBART BROTT MOT PAKTEN Gå försiktigt . 
Patrick Kennedy . 
Stå stilla . 
Ett bra råd . 
Det känns inget vidare när jag gör det . 
Om ni kommer närmare kastar jag mig ner i hålet . 
Vi stannar här , men ditt sår behöver behandlas . 
Alltså , det är lustigt , det verkar som om ni kommer att ge mig nya sår med era vapen . 
Du är en rymling som sågs brandbomba min station . 
Du förstår varför vi är lite försiktiga . 
Vi kan hjälpa dig . 
Jag litar inte på er . 
Det är därför jag är här i mörkret och blöder i ett jävla hål ! Vi har första hjälpen - i generatorrummet . 
Väntade du på det ? 
Skjuter du mig nu när vi är ensamma , och hoppas att vicesheriff Långhårig inte räknade skotthålen ? 
Vi skjuter inte folk som inte utgör ett direkt hot . 
Jag utgör ett direkt hot . 
Med allt jag vet , vore det bäst för dig att gå . 
Det kan jag inte göra . Jag svor en ed . Där ingår att vårda skadade . 
Vårda skadade ? 
Inser du inte att allt är lögn ? 
Allt de sa åt oss . Pakten . Den är för att hålla oss i schack . Och vi får aldrig veta sanningen . 
Hellre skulle Sims skjuta oss allihop . 
Känner du mr Sims ? 
Ja , jag känner honom . 
Jag hjälpte Nichols . 
Jag greps och förhördes . Varför tror du att jag är här nere ? Berätta . Okej . Jag ska berätta . 
Ge mig pistolen , bara . 
Just det . Du kan inte , för du litar inte på mig . 
Om du ska skjuta mig , ber jag dig att skjuta mig i pannan . 
Snälla . 
Jag hittade det här i Juliette Nichols lägenhet . Inuti en bok . 
Jag förstörde resten . 
Jag vet inte varför jag sparade det . 
Om du berättar för nån om det , är jag rökt . 
Skaffa hit en läkare . Inte en vicesheriff med plåster . Då ska jag berätta allt du vill veta . Nej , jag ska berätta allt du säkert som fan inte vill veta . 
Nya villkor . 
Hur lång är kabeln ? Det lär du märka . 
Den här ? Den är inte Juliettes . Så förbanne mig om jag låter dig sälja den som hennes . 
Barnes , stanna inte . 
Kom . 
- Nån uppdatering ? - Inte än . Sök efter två personer som rör sig nedför trappan . Uppfattat . 
Nivå 92 . Två bärare på väg ner . 
Jag är strax bakom . Meddela borgmästaren . 
Uppfattat . 
Här är mat . Vad gör du ? 
Jag försökte spåra upp en hjälm som stals från dräktrummet . 
Så jag gick till en anställds lägenhet för att hitta den . 
Trina Samuels lägenhet . 
Trina Samuel . 
Ja . Hon var Solos flickvän . 
Ja . Jag har inte tänkt på henne på länge . 
Faktiskt tycker jag inte om att tänka på henne . 
Vill du ha kyckling eller nötkött ? 
Varför ljuger du för mig ? 
Jag vet inte vad du menar . 
Solo , Trina . Det där är hon . Men det där är inte du . 
Nej . För ... Titta . Jag hittade det här . Cole Myers , IT-skuggan . 
- Det är den verkliga ... 
- Jag är IT-skuggan ! 
Du vet inte vad du pratar om ! 
Säg inte de där orden till mig ! Aldrig nånsin ! 
Jag är Solo ! 
Jag är IT-skuggan , hör du det ? 
- Okej . 
- Jag är Solo ! Jag är IT-skuggan ! Du är Solo . 
Du är Solo . 
Förlåt mig . 
Förlåt mig . 
Du ser bedrövlig ut . Du borde äta nåt . 
Jag är inte hungrig . 
Jag mår inte bra . 
Jag behöver ... Jag ska gå och lägga mig . 
Jag ska bara ... Är det tillräckligt långt ner ? 
Jag tror det . 
Men kommer det att hålla för din tyngd ? Det vet jag inte . 
Mekaniska ! 
Stanna ! 
- Helvete . - Fan . 
Kom igen . 
Det finns ingen broms , va ? 
Vi har kabeln , och så slutet på kabeln . 
Vi dör åtminstone på Botten . 
Ge mig din hand ! 
Se upp . 
- Där är de ! 
- Ta dem ! 
Se upp ! 
- Helvete ! - De kom igenom , sir . 
Jag märkte det . 
Håll den här kanalen öppen . 
Sheriff Billings , hör du mig ? 
Sheriff Billings . Ja , borgmästaren ? Jag måste tyvärr meddela att rymlingarna från Mekaniska just blev ditt problem . 
Som Silons lojala tjänare vet jag att du kommer att gripa dem . 
Självklart , borgmästaren . 
Du vet att jag alltid kommer att troget tjäna Silon och Pakten . 
Kom igen . 
