Patrull V7 från inspektör Lenker . Jag går in i Hatherways Flats , nionde våningen . Jag går mot lägenhet 942 , misstänkt på fri fot . 
- Lenker , patrull 7 , uppfattat . 
- Gå in . Vi är på väg . Framme om tre minuter . Fortsätt med försiktighet . 
Polis ! 
- Går in . - Uppfattat . Kommer om två minuter . 
Nej , stanna ! 
Polis ! 
Stanna ! 
Han är det . 
" Clive Silcox . " Det är absolut han . 
Han finns i databasen , vad har han gjort ? 
Ett antal anmälningar , misshandel , våld i hemmet , medlem i en förbjuden organisation . Nån ultrahöger , Combat League tror jag . 
Inget som ledde till fällande dom . 
Hur långt tillbaka går anmälningarna om misshandel ? 
Augusti 2009 . 
Polisen kallad till bråk på Michaels Street . Michaels Street . Han bor lokalt . Varför är det intressant ? 
Offret , Maria De Souza . 
Jag tror att hon var uppringaren från Hayes Lane i tisdags kväll . 
Det anonyma larmsamtalet ? Ja , sir . 
Våldsam pojkvän som hävdat att han dödade Adelaide Burrowes . 
Jag begärde förstärkning , om du minns . - June ... - Och nu ... Han kan ha grannar , vänner från jobbet , ex-partners . 
- Om han har en historia av tvång ... - Hör på ... Nej , jag hade honom . 
Du gjorde ditt bästa . 
Det viktigaste är att du är okej . 
Det är det viktiga . 
Så här , om det är nåt skumt med det här andra mordet , Adelaide Burrowes ska vi utreda det . 
Oavsett vem som felat . 
Ju större de är ... Kim . Vad kan jag göra för dig ? ... desto hårdare faller de . 
Bri . Jag hörde att du har ett mord i ditt distrikt . 
Ursäkta mig . Hej . Jag söker June Lenker . 
- Hon kom in hit för ett tag sen . - Helvete . 
- Mår du bra ? - Jadå . 
- Säkert ? - Ja . 
Kom . 
Vad har de gjort med dina kläder ? 
De tog dem för att kolla fibrer och DNA ... - Det är normalt . - Jaha . Normalt ? Det finns inget normal med det här . 
Leo , det är ingen fara . Bara jack och skråmor . 
Förlåt , jag vet inte vad det är med mig . Det är okej . Bara ... vänta lite . 
Ursäkta mig . Ursäkta . Allt är bra , vännen . Finns det nån läkare här ? För min fru är polis och har blivit misshandlad . 
Leo . Leo , jag har klartecken att gå hem . 
Jag väntar bara på att läkaren ska skriva ut mig . Hon behöver träffa en läkare . - Okej ? - Okej . - Får hon träffa honom nu , tack ? - Ett ögonblick . Tack . 
Det är okej . Det är okej . 
Raring , vad gör du ? Inget . 
Är det vad jag tror ? 
- Lägger du ut det på sociala medier ? - Nej . 
Jösses , det gör du . Får jag se . 
- Kom igen , mamma . - Oj , alltså . Jacob . Alltså , vad gör du ? Du lägger ut din mammas skador på nätet . Hoppas att din pappa inte följer dig . 
Nej . Jag har blockerat honom . 
Men jag har fått 13 gilla och det ökar . Är det bra ? 
Du låter typ 80 år gammal . 
Nån kallade mig just en tuffing . 
Det kan jag leva med , " tuffing " . Förlåt . 
Är det vad som krävs för att du ska vara stolt över mig ? 
Det är han . 
Clive Silcox . 
Det här är Clive Silcox . 
Så , alla som kan ha råkat på honom . Ex-flickvän , syster , familj . 
Allt hjälper . 
STOPPA VÅLD I HEMMET Och det här är mitt direktnummer . 
Det här är mitt nya nummer . 
Tack , raring . Precis vad jag behövde . Mjölk , en sockerbit ? 
Två , faktiskt . Det går utför . 
Nej , ingen fara . Tänk att du jobbar kväll än ? Man vänjer sig . 
Jag lägger inte ner min själ i det . Det är bara jobb . Det är en chansning , men jag försöker spåra upp en man , Clive Silcox . 
Jag ska fråga runt . 
June , det har hänt saker i fallet Hatherway Towers . Ring mig är du snäll . 
Ursäkta mig . 
Sir . Vet du att jag var först på platsen ? 
Låt mig stoppa dig där . 
Det visar sig att den här Silcox redan är föremål för en utredning . Verkligen ? Ja . Tydligen en ung kvinna som överfölls på väg hem i oktober . 
Samordnarna ansåg det bättre att existerande team utredde det här mordet . 
Har ni hittat honom än ? 
Jag hänvisar alla frågor till min kollega , inspektör Gearing . 
Hon gör jobbet , jag är bara här för syns skull . 
Vänta , så ... Tror hon att han är kvar här ? 
Det där ser inte bra ut . 
Sir , innan offret dog , Maria , identifierade hon sig för larmcentralen som uppringaren från Hayes Lane . 
- Uppringaren från Hayes Lane ? - Det anonyma samtalet ... - ... jag visade dig i onsdags . - Visst , ja . Så om ni lyckas gripa den misstänkte , ber jag om tillstånd att förhöra honom om anklagelserna . 
- Anklagelser ? 
- Mordet på Adelaide Burrowes . 
Två samtal , samma kvinna . Är det din hypotes ? - Ja . 
- Mycket tunt . 
Nej . Maria De Souza ... Hon sa till telefonisten : " Vi har pratat förut ... " 
Ja , pratat förut . Hon sa inte var . Hon sa inte när . 
Vi kan inte bara ignorera det . 
Det finns fysiska likheter mellan kvinnorna . 
De har samma kroppsbyggnad . De är båda spansktalande . De låter likadant . 
De sa att du såg henne falla . 
Ja . Jag vill inte förefalla överlägsen , men jag hörde en inspelning av samtalet och vad du sa . Rådet du gav de sista ögonblicken i hennes liv . Det var helt rätt . Du gjorde rätt . Du var hos henne . 
Hon var uppringaren . 
- Okej . - Hon är uppringaren från Hayes Lane . 
- Och det är troligt ... - Man ser vad man vill se . Så gör vi alla . 
Jag vill bara förhöra mannen . 
Samma här . Men tyvärr har vi inte hittat honom . 
Det har gått tio timmar . Ni slösar bort tiden . 
Jag tillskriver det där din bula i huvudet . 
Jag mår bra . Nej . Du var offer för en misshandel . 
- Varför tror ni att han är kvar ? 
- Det är ingen baksmälla . 
Ni slösar tid och resurser . - Ni borde vara ute och leta . 
- Gå hem . Få lite sömn . 
Vi är på samma sida . 
Hör på . Han hade en flickvän för länge sen . 
Hon var som jag . 
Han sa : " Dumma slyna . Hon lyssnade aldrig . " 
Hon gjorde honom aldrig nöjd . 
- Kan du säga ditt namn ? 
- Maria . 
Okej , Maria . 
Jag ringde . Jag pratade med dig tidigare . 
Ja , jag minns . 
Han högg henne många gånger med samma kniv som han högg mig . 
En man har fått 24 års fängelse för mordet på henne . Han säger att den här killen i Whitecross ... Han säger att han är en nolla och en ... Din dumma slyna . 
- Säg att du förstår . 
- Få tag i henne ... - " Dumma slyna . Hon lyssnade aldrig . " 
Hon gjorde honom aldrig nöjd . 
Vi har gjort en lista över dina fordonssökningar i databasen . 
Som du ser finns inget aktnummer för nån av dem . Inget brott . 
Så vi vill att du går tillbaka till varje sökning och lägger till det relevanta aktnumret . 
Som du säkert vet bryter det mot ... Gå tillbaka i din arbetslogg , gräv fram aktnumren och ordna till det här . 
Sir , jag vill göra en röstanalys på de två nödsamtalen . Hayes Lane och gårdagens offer , för att bekräfta om det är samma kvinna eller inte . 
Det är inte vårt fall , June . Det har klargjorts . Sir . Uppringaren från Hayes Lane anmäldes av kontrollcentret . Du bad mig följa upp det . 
Om uppringaren var Maria De Souza kan vi avsluta fallet . Det är allt . Okej , hör på . 
Jag ser att du är upprörd . Okej . 
Men tänk lite på Jim . Han saknar folk till inbrotten i Oakmoor . Visst ? - Ja , sir . - Så du kan väl jobba med det ? 
- Allt kommer att ordna sig för dig . 
- Jag vill inte att folk ska glo . 
Kom igen . Du är bruden , raring . Det är din stora dag . Du måste visa upp dig . 
Är du Doris Mathis ? Ja. vi är nästan klara här . Gå in , bara . 
Jag vet inte . Kom och titta i spegeln . 
- Oj . - Ja , du ser ? 
- Vi ses nästa vecka . - Okej . Vi ses då . 
- Hur kan jag hjälpa dig ? - Hon blir jättefin . 
Åh , tack . 
Jag är kriminalinspektör June Lenker . Ursäkta att jag stör . Okej . 
Latisha , ursäktar du oss ett tag ? Visst . 
Vi försöker spåra den här mannen . 
Han heter Clive Silcox . Han är efterlyst . Vi försöker ta reda på var han gömmer sig . Han bor i trakten . 
Så vi kontaktar alla som kan ha råkat på honom eller kan ha varit bekant med honom . 
- Så , kanske du ... - Säg mig , vad gör en rar kvinna som du i polisväsendet ? 
Kanske din son ? De kanske kände varandra förr . 
Har du pratat med min Errol ? Nej , hur så ? Tror du ... Tror du att de kände varandra ? 
Han kanske var hemma hos Errol ? Han kanske kände Adelaide ? 
Adelaide ? Varför nämner du henne ? 
Hör på . Jag är ingen novis . Jag kan genomskåda skitsnack . 
Jag försöker bara få lite hjälp . 
Har du legitimation , ms ... Vad var det ? 
Lenker . June Lenker . 
Lyssna noga på mig , inspektör Lenker . Om du tror att du kan valsa in här och försöka sätta dit min Errol för nåt nytt ... - Det är inte det jag försöker göra . - Gå härifrån . 
Vem skickade dig ? 
Skickade han dig ? - Vem då ? 
- Hegarty . 
Och hans gäng . 
Hans gäng , de bara ljuger . Och de ... De burade in min son , vet du . Och när man försöker stå där artigt och säga : " Ursäkta , ni har nog gjort ett misstag här . " Ett misstag ! Bara det . 
Hälsa honom från mig : " Jag är fortfarande här . " 
Okej . Clive Silcox . 
I mars 2011 bodde han på 24B Lake Street . 
Lake Street . Här i närheten . 
Anställd hos Rudin ' s. Leveranser . 
Det gamla yiddish-stället ? 
Nåt alibi ? 
Inte vad jag kunde hitta . 
Synd . Och vi förhörde honom aldrig då ? 
Självklart inte . 
Vadå ? Vi kan väl inte förhöra varenda skummis i London ? 
Nä , vi hade gripit vår man . 
Hör på , allt som placerar Silcox nära Adelaide , Errol Mathis eller våningen ... Allt hon kan använda mot mig eller utredningen , vill jag ha reda på . Okej ? 
Jag trakasserade henne inte . Men så upplevde hon det . 
Så berätta för mig vad min klient har att göra med Clive Silcox , annars anmäler jag dig för tjänstefel . 
Det är möjligt att Silcox har information som är relevant för mordet på Adelaide . 
Så allt som kopplar Silcox till Adelaide eller Errol ... 
" Relevant information " ? Vad menar du ? Var han ett vittne ? Eller en misstänkt ? 
Jag kan inte ... Det är konfidentiellt . För Guds skull . 
- Chloe ? 
- Ja ? Du har kompisar i Hackney Downs , va ? Ja ? 
Jag behöver en tjänst . Alltså , om det gäller ditt mordfall ... - Kom igen , Chloe . - Jag vägrar bli inblandad . 
Jag kan inte lägga mig i . Det är konfidentiellt . Snälla . Jag skulle inte be dig om det inte var viktigt . 
Hur stor är tjänsten ? 
- Varsågod . - Tack . 
Starkaste kaffet i Dalston . Tacka inte förrän du har smakat . 
I alla fall , jag pratade med Doris , och Errol gick i skolan med honom . 
- Med vem ? 
- Clive Silcox . 
St . Joseph ' s Academy . 
Men Clive var typ två år äldre , så de var inte kompisar direkt . Men Doris kände familjen , sa hon . Lite grann . Lite grann ? Hur då ? 
Errol hade en kusin , Jameel , som var förtjust i Silcox syster . Men Doris satte ner foten , så ... Så Errol kände honom ? Det gjorde han . 
Tack . 
Ingen orsak . 
Tycker du att jag har en aggressiv framtoning ? 
Aggressiv ? Till exempel ? Till exempel rastlös . 
Enveten . Dominerande . Tokig . Lägg gärna till nåt om du vill . 
Roy sa att jag var upprörd . Men det är ju bara omskrivning för galen kärring , eller hur ? 
- June ? 
- Vadå ? 
Du har genomgått ett trauma . Han har rätt att fråga . 
Så jag övertänker . 
Du parkerar sexigt , vet du det ? 
En märkligt nischad komplimang . 
Så där ? 
- Så där ? - För fan . - Vill du göra färdigt själv ? - Nej . Jag kan gå och köpa glass så länge . 
Känner du dig stabil ? 
Jag sitter i en knipa , faktiskt . 
Heja . 
Passa , passa ! 
Jag fattar inte . Så du sökte i en databas , än sen ? 
Alla sökningar måste vara jobbrelaterade . Man ska bifoga ett aktnummer . 
Och ? 
Det var inte för mig , utan för mamma . 
Okej , hur många gånger ? 
Vet inte . Åtta ? 
Åtta ? June . 
Varför sa du inget ? 
Jag visste vad du skulle säga . Och jag vill inte att hon blir intagen igen . Det får inte hända . Aldrig mer . 
Så det är lösningen ? Att göra illegala datasökningar ? Inget av det här hade hänt om det inte var för den där jäveln . - Hegarty . Bla-bla . - Du blev slumpvis kollad , sa du ju . 
Han har inflytande . Han känner folk . Okej , stäm i bäcken . Prata med din chef . 
- Roy ? 
- Berätta vad du gjorde , stor sak . 
Det är bokstavligen det värsta jag kan göra . 
- Varför ? - Han är samvetsgrann och känner sig tvungen att rapportera det . 
Okej . Gå högre upp i näringskedjan . Prata med vice polischefen . Han du pratade om , som ville ha dig som kriminalinspektör . 
Jaha , bara ringa upp honom ? " Hej , minns du mig ? 
Jag är kvinnan du var trevlig mot vid en rekryteringshelg i Hounslow . " - Varför inte ? 
- För jag är inte du . 
Jag går inte genom livet och tar mig själv för given . 
Det är inget fel att vara självsäker . Självsäker ? 
Jag är inte helt säker på vad det betyder . 
Jaha . Så det handlar om vitas privilegier . Jag vet inte , Leo . 
Men jag vet att jag inte skulle skälla på nån stackars akutsköterska bara för att jag har lust att avreagera mig . 
- Är man självsäker då ? Jag vet inte . Kanske . Troligen . Jag vet inte . 
Vad pågår ? 
- Han fällde honom . - Gjorde han ? 
Ja . Krokben . 
Jake , lyssna på domaren . 
Du får en varning nu . En gång till så blir du utvisad . Okej ? Okej . Spela på . 
Kom igen , Jakey . Upp med hakan . 
Hör på . Jag ber om ursäkt om jag var oförskämd mot en sköterska , men jag var uppriven . 
Jag var upprörd för att jag just hade fått ett samtal . 
Och ett tag ... Lyssnar du ens ? 
Jag trodde att du var död . 
Kom igen , kompis . 
Vet du ibland vet jag inte om vi befinner oss på samma planet . 
Det här är Becca från härbärget på Moore Street . 
- Ja . Hej . - Du frågade om Clive Silcox ? 
- J ? - Vi har funnit ... Det är jobbet . 
Jaha , då tar vi väl bussen , då ? 
Nån har trätt fram ... Okej . Inga problem . 
Hej , är du Dawn ? Dawn Taylor ? 
- Det stämmer . - Ursäkta att jag stör . Jag är kriminalinspektör June Lenker . 
Jag försöker hitta en man som du kände tidigare , Clive Silcox ? 
Ni kände visst varandra 2018 . 
Har du nån aning om var han kan finnas ? Eller några vänner ? Platser där han kan ... 
Följ med mig . 
Okej . Tack för din tid . Varför inte ? Min mamma . 
Zero Yankee Delta . Det här är inspektör June Lenker . 
Jag är på Verlaine Road 70 . 
Jag tror att jag har hittat Clive Silcox . 
Uppfattat . 
Understöd är på väg . 
Hur långt bort ? Zero , delta , bravo . Framme om sex minuter . Sex minuter bort . Stanna där du är . Vänta på förstärkningen , kom . 
Uppfattat . 
Zero Delta Yankee . Det är bråk inne i huset , kom . 
Avvakta . Förstärkning är på väg . 
Så fan heller . 
Polis ! Öppna dörren . 
Polis ! 
Zero Delta Yankee . Det pågår misshandel inne i huset . 
- Vad händer ? 
- Får jag använda din trädgård ? - Jadå . - Avvakta förstärkningen . 
Zero Delta Yankee . Skicka brandkår genast . 
Zero Delta Yankee , upprepa . 
Zero Delta Yankee , upprepa . 
Zero Delta Yankee , upprepa . 
Jag sa att huset brinner ! 
Skicka brandkår genast . 
Dawn ? 
- Är det nån här ? - Hjälp ! 
Vi är här inne ! 
Undan från dörren ! 
Ut ! Nedför trappan ! Fort ! 
Det här kom inte från mig . 
Svär . 
Har du patolograpporten ? Svär . 
Jag svär . 
Radera den så fort du är klar . Ja . 
Redo ? Jadå . 
Vet han att jag kommer att sitta med ? Ja . Han föreslog det faktiskt . 
Tack båda två för att ni tog er tid ... - Det är det minsta vi kan göra . - Så , senaste nytt . 
Clive Silcox har erkänt mordet . Fantastiskt . 
Han erkände utan omsvep . 
Mordet på Maria De Souza . Våldsamt motstånd mot polis . 
Han gav sig på fel polis den här gången . Verkligen . 
Vi frågade : " Varför dödade du henne ? " Han sa : 
Hon spillde färg på mattan . - Nej . - Färg på mattan . 
När man tror sig ha hört allt . 
Åklagarämbetet gav klartecken , vi åtalade honom för tre timmar sen . Så allt är klart . 
Jag vill ha tillstånd att förhöra Silcox . 
- Angående ? 
- Mordet på Adelaide Burrowes . 
Det är ett gammalt fall . Det var ... 2011 . Det är ett gammalt mord . 
Pojkvännen , Errol Mathis , avtjänar ... - Tjugofyra år . - Ja . Jag vill bara prata med honom . 
Jaha . Okej , jag tycker att vi ska rensa luften här . Och hitta en lösning . 
Inspektör Le ... Får jag kalla dig June ? 
- Visst . - Okej , June . 
Vilken ny information har du som placerar Clive Silcox i lägenheten med Adelaide Burrowes ? 
Han bodde i trakten då . 
24B Lake Street . Det stämmer . 
- Bara 500 meter från Towers . 
- Det stora gamla kvarteret . 
Silcox har en historia av anklagelser för våld mot kvinnor . En gång 2009 , och sen ... Maj 2011 . Ja . Vad mer ? 
De gick i skolan ihop . Silcox och Errol Mathis . 
St . Joseph ' s. Över 2 000 elever . 
Flera års åldersskillnad . 
Silcox hade en syster , Leanne , som var kompis med Errols kusin . Kusin ? Vi har alla kusiner . En del fler än andra . 
Pratade ni ens med honom ? - June ... - För att avföra honom från utredningen ? 
June , känner du till uttrycket " omedveten bias " ? 
Jag gick kursen . Fick diplomet . Det var väldigt lärorikt . 
Du förstår , grejen med omedveten bias är ... Jag vet vad omedveten bias är . 
Nå , jag förklarar för de tröga . Ursäkta , Roy . 
Du vet , ibland kan en polis ha en förvrängd inställning till ett fall . På grund av sina , ursäkta mig , redan existerande fördomar . Fördomar . Fördomar ? 
Okej , vi möts på halva vägen . Tro ? 
Övertygelse ? Är det okej ? 
June här har en övertygelse om att denne Errol Mathis , en man av västafrikanskt ursprung har blivit orätt dömd av skäl som är dunkla . Fast det kom ett nödsamtal . 
Försök igen . Två samtal . Två kvinnor . 
Två samtal . En kvinna . 
Vi kan inte ... Vi kan inte utesluta det . 
Vet du hur många kvinnor som utsattes för våld i hemmet i den här stan bara i fjol ? Visst vet du det . 
- Nästan en kvarts miljon . - Ja . Nästan en kvarts miljon . 
Båda var portugisisktalande . Det är många som talar portugisiska . Vi pratar om 80 000 eller 90 000 . 
Och därför bör vi utföra röstanalys ... Men för jösse namn . ... för att bekräfta om det var samma kvinna som ringde , eller inte . Okej . 
Hon då ? Maria ? 
Vem ? Jo , offret . För att inte tala om labbkostnaden . Vi har femsiffriga budgetöverdrag . 
Vi har en man i häkte som är villig att erkänna mordet på henne . 
Vilket besparar hennes mor , bror och två moderlösa pojkar en jobbig rättegång . 
Hennes kropp är redan på väg hem till São Paulo . Det är goda nyheter . Men du vill riva upp alltihop på grund av din käpphäst . 
Maria hade två gamla knivsår . 
Axeln . Buken . 
Uppringaren från Hayes Lane sa också att hon hade knivhuggits av sin partner . Och hon sa : " Han knivhögg henne " , alltså Adelaide , " många gånger med samma kniv han högg mig . " 
Ursäkta , varifrån kommer det här ? 
- Hennes ord från telefonsamtalet . - Jag menar inte det . Jag menar ms De Souzas skador . 
June , har du sett patologirapporten ? 
Det viktiga här är ... Nej . Förlåt att jag tjatar , men patolograpporten sändes väl konfidentiellt till Viv och hennes team ? 
Ja ? Så om inte ... Viv , delade du den med inspektör Lenker ? 
- Nej , sir . - " Nej , sir . " 
Så jag måste fråga , hur hamnade den på ditt skrivbord ? 
Delade nån den med dig ? Nej . 
Så vadå ? Är du en hacker i maskopi med Nordkorea ? 
Påstår du att du inte har läst patolograpporten ? 
Nej , sir . 
Så var fick du informationen ? 
Jag såg dem . 
Du såg dem ? 
Jag var först på platsen . 
När jag fann Maria kollade jag givetvis hennes livstecken . Jag såg dem . 
Jag såg hennes skador . 
Två gamla skador . På en sekund . 
Två uppringare . Matchande knivsår . 
Är det verkligen en slump ? 
Kör . 
Ren mottagning . Allt handlar om timing . Man måste ... Du ser ? 
Ja ! Jättebra . 
- En gång till . - Okej . 
Kom igen , tackla mig . 
Vad är det här ? Extra träning ? Okej . Kom igen då . Vänta lite . Vänta . Okej . Vänta . 
Vilket mål ! 
Du lär dig allting av mig . - Allting av mig . - Mamma , det är hands . 
Du skämmer ut dig . 
En gång till . 
Du fick som du ville . 
Med tanke på " de exceptionella omständigheterna " . 
Fången kommer ut . 
Du har klartecken att prata med den misstänkte . Tack . 
Men dina frågor gås igenom i förväg , okej ? Okej . 
Specifika referenser till mordet på Burrowes är förbjudna . Förstått ? 
Okej . 
Annars är det bara att köra . 
Tack , sir . 
Clive Silcox , du har erkänt mordet på Maria De Souza . Men jag är här för att fråga dig om en annan sak . 
I mars 2011 bodde du på 24B Lake Street . Stämmer det ? 
Känner du igen den här mannen ? 
Känner du honom ? 
Errol . Errol Mathis . Ni gick på St . Joseph ' s samtidigt ? 
Kände du familjen ? Roy . 
Är du medveten om att Errol Mathis - avtjänar ett långt fängelsestraff ? - Tack . 
Tjugofyra år , va ? Stämmer . Vet du var ? 
- Whitecross ? 
- Whitecross Prison , det stämmer . 
- Än sen ? 
- Inspektör Lenker . 
Vet du varför ? Ja . - Ursäkta ... - Det är allmänt känt . Om du försöker snärja min klient ... Nej . Jag vill bara att han säger det . 
Vad heter hon ? 
- Okej . - Säg det . 
Säg hennes namn . 
Jag avslutar den här intervjun . Klockan är 14 : 36 . 
Vad fan snackar hon om ? 
- Han kände dem . Han kände dem båda . - June . 
- Dan , vill du ... - Nej . Gör det du . 
Med tanke på din begäran ansåg Hegarty det klokt att villfara den och köra en röstanalys på de två nödsamtalen . 
Den är definitiv . 
Fonetikern och teknikern nådde samma slutsats . Olike betoningar . Olika vokalljud . Två olika kvinnor . - Va ? 
- Det är utom allt tvivel . Uppringaren från Hayes Lane var inte Maria De Souza . 
Inget överhuvudtaget binder Clive Silcox till det gamla mordet . Ja ? 
Är vi överens ? Låt oss avsluta det här en gång för alla . 
Okej ? 
Vad är det med dig ? 
Se på Chloe . 
Hon har inga problem . 
Hon bara sköter jobbet . 
Och granskningsgruppen ? Har du hört av dig till dem ? Inte ? 
Se till att göra det . Annars anmäls du för tjänstefel . 
Han hade rätt . Jag hade fel . 
Helvete . Jag avskyr sånt . 
Hör på ... Det går ett rykte . 
Dagen efter att Silcox mördade Maria De Souza fick Hegarty röstanalysen gjord på direkten . 
Va ? 
Han visste att det var två uppringare och ... Han satt på rapporten . 
Vänta . Hela det där mötet . Ge klartecken till intervjun . Varför ? Varför gjorde han det ? 
Man måste exploatera situationen . 
Han lurade mig . 
Det var en fälla , och jag gick rakt i den . 
Han vill trycka ner mig i skoskaften så att jag håller tyst sen . 
Inte jag . 
Han hade en flickvän för länge sen . 
Han sa : " Dumma slyna . Hon lyssnar aldrig . " Hon gjorde honom aldrig nöjd . 
Han högg henne många gånger med samma kniv som han högg mig . 
En man har fått 24 års fängelse för mordet på henne . Och han säger att den här killen i Whitecross ... Han säger att han är en sån nolla och ... När hände det här ? 
I tisdags . 
De här samtalen är konfidentiella . 
Om du berättar för nån , kommer de att krossa mig . 
Här . 
Jag trodde att du var muslim . 
Jag är sikh , du vet . Singh ? Sonya Singh ? 
Vi dricker sånt här som Lucozade . 
Okej . Du hade fel . 
Du förlorade kampen , bu-hu . Men vet du vad ? Hon är vid liv . 
Hon är den enda som kan hjälpa Errol , och hon är vid liv . 
Ja . Och vi ska hitta henne . 
