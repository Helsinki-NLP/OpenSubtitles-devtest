Det är vad alla kallar mig , som ett tecken på kärlek och respekt . 
Samsik eller farbror Samsik . 
Jag älskar det . Jag älskar mitt smeknamn . 
När den är byggd blir jag officiell medlem i Cheongwooförbundet . 
Vet du vad det betyder ? 
Jag blir den som störtar adeln . 
Vi äntligen äta pizza som amerikanerna . 
Ni har nog aldrig hört talas om pizza . 
Det är jättegott . 
Rekonstruktionsbyråns chef , Kim San . 
Han studerade ekonomi i USA med ett Albrightstipendium . 
Herrn . 
Yoon Palbong från Dongdaemunligan . 
Vill du ha hans område ? 
Yoon Palbong skickar 25 män till Innovationspartiets tal . För att föra liv under herr Choo Intaes tal . 
Yoon Palbong får inte komma undan . 
Se till att bryta hans ben , okej ? 
Jag ska lära honom en läxa på Innovationspartiets tal . Oroa dig inte . 
Döda Yoon Palbong . 
Ursäkta ? 
I USA var allt överflödigt och vackert . Men mitt land var slitet och mitt folk svalt . 
Vet nån vad pizza är ? 
Du vet hur pizza smakar . 
Har du verkligen smakat det ? 
Seohae Olja , Sail Utveckling Vd Pak Doochill 
Jag ser i folks ögon om de har vad som krävs . Frågar du mig , kan du bli president en dag . Men låt oss vara ödmjuka och säga minister . 
Ska jag kalla dig minister ? 
När kan det implementeras ? 
Jag kan ge dig ett tydligt svar . 
Gör slut med Choo Yeojin . 
Du kan inte förverkliga din dröm som Choo Intaes svärson . 
Rekonstruktionsbyrån ska läggas ner . 
Jag ger inte upp rekonstruktionsprojektet . 
Har du lämnat inrikesministeriet ? 
Finns det en plats i Innovationspartiet ? 
Vårt parti är inte redo än . 
Hur mycket jag än försöker , kan jag inget göra . 
Varför skakar du inte om denna obevekliga värld ? 
Jag har en dröm . 
Jag vill förändra vårt land till det bättre . 
Det är ingen dröm . 
Det är hyckleri . 
Hyckleri förklätt till en dröm . 
Lägg då all din uppmärksamhet på det du vill uppnå ! 
Jag vill göra det ! 
Jag vill genomföra nationella rekonstruktionsprojektet ! 
Jag gör slut med henne . 
Gå bara . 
Allt man vill ha i livet har ett pris . 
Jag har en storslagen plan för hur Cheongwooförbundet ska ta över landet . 
En storslagen plan ? 
Vi inför ett parlamentariskt system och mutar hela nationalförsamlingen . 
Måste vi döda Yoon Palbong direkt ? 
Han behövs i nästa val . 
Nej . 
Låt Taemin ta hand om honom . 
Han hyser nog agg mot Yoon Palbong . 
Vem vill han se död nu ? 
Döda honom , så kan du börja om i Osaka . 
Jag har bevis på Kang Seongmins inblandning i Sineuialliansen . 
Kang Seongmin vill att jag dödar dig . 
Jag är här för att rädda dig . 
- Flytta på dig , jävel . 
- Du din ... 
Hördu , Haejun ! 
Fan ! 
Haejun ! 
Kang Seongmins far dog i en explosionsolycka . 
Sineuialliansen var kända för sina bomber . 
Enligt polisrapporten sköts Yoon Palbong först . 
Han var inte ute efter Choo . 
Uncle Samsik 
Uncle Samsik 
Hallå ? 
Minister Kim . 
Hej . 
Välkommen . 
Varför ville du träffas så sent ? 
Känner du Cha Taemin från Sineuialliansen ? 
Va ? 
Presenterade du Yoon Palbong för Kwangmin med Innovationspartiet i åtanke ? 
Ja . 
Tipsade du media om Kang Seongmin ? Ja . 
Varför då ? 
Jag tar kaffet sen . 
Yoon Palbong utförde mycket skitjobb åt Kang Seongmin . 
Det gjorde jag också . Men Yoon Palbong förrådde Kang Seongmin . 
- En kaffe , tack . 
- Okej . 
Hur förrådde han honom ? 
Jag kan inte berätta detaljerna . 
Du vill jobba för vår gemensamma dröm . Hur kan vi jobba ihop med alla hemligheter ? 
Det är bäst om du inte vet . 
Angående herr Choo ... 
Beordrade du hans mord ? 
Du låter fantasin flöda igen . 
Jag gjorde slut med Yeojin . 
Vad har du gjort under tiden ? 
Du har hemligheter och smider farliga planer i smyg . Men jag ska stå på din sida ? 
Du läste väl artikeln om ledamot An Minchul , An Yosubs son ? 
Yoon Palbong och jag dödade honom . 
Tre år tidigare 
Säg till om ni behöver hjälp i distriktet . 
Så generöst av dig . 
Vi är dig evigt tacksam . 
Ledamot Kang . 
Trevligt . 
Du ville ses ? 
Säkerhetschefen sa nåt intressant när vi tog en drink . 
Vad sa han ? 
Cha Taemin från Sineuialliansen . 
Du växte väl upp med honom ? 
Anarki , knappast . 
De har dödat dina rivaler . 
Smart drag . 
Låt mig låna Sineuialliansen nån gång . 
Vi måste dela med oss . 
An Minchul har avslöjat oss . 
Seongmin . Du borde sluta nu . 
Vad menar du ? 
Jag åker till Osaka med de andra . 
Farbror Samsik kan fixa jobb . 
Jag tror inte att jag klarar detta . 
Var inte sån . 
Jag räknar med dig . 
Cha Taemin lydde inte Kang Seongmins order . 
Herrn . 
Den här mannen erkände på vägen tillbaka . 
Kan du ta fast Chae Taemin ? 
Visst , mina män hämtar honom . 
Varför släpper du inte Taemin ? 
Det här är killen som hanterade bomberna i alliansen . 
Låt mig ta honom och sen tar vi itu med An Minchul själva . 
Det låter bra . 
Kan du hjälpa oss lite mer , herr Yoon ? 
Gärna . 
Vad vill du ha i gengäld ? 
Min dröm är att bära nationalförsamlingens emblem . 
Nominera mig till Dongdaemun , så gör jag vad som helst . 
Det finns en jävel . 
Kang Seongmin beordrade Yoon Palbong att hämta Cha Taemin . 
Skulle du komma undan helskinnad ? 
Säg till Kang Seongmin att jag inte ställer upp mer . 
Era förrädare . 
Trodde ni att ni kunde gömma er utan att åka fast ? 
Ni kan rädda er själva . 
Det är enkelt . 
Ska jag slänga er i havet eller låta er jobba ? 
Jag jobbar för dig . 
Jag också . 
Jag med . 
Han drömde om en plats i nationalförsamlingen , så Yoon Palbong ställde upp . 
Han fångade Taemin innan han dödade An Minchul . 
Minchul ! 
Cha Taemin förrådde Kang Seongmin , så Yoon Palbong och jag dödade An Minchul i hans ställe . 
Yoon Palbong tjatade om det , så vi dödade honom . 
Varför visa honom Innovationspartiet ? 
Han var besatt av nationalförsamlingen , så jag trodde att en nominering skulle tysta honom . 
Nyhetsartikeln , då ? 
Den skulle ruinera Kang Seongmin . Han är ett hot . 
Vi måste gradvis försvaga hans makt för att störta honom . 
Var är Cha Taemin nu ? 
Han gömmer sig . 
Herr Cha . 
Herr Cha ? 
Vänta , det finns en dörr här . 
Rör dig inte . Vem är du ? 
Var är Cha Taemin ? 
Jag letar efter honom . 
Du är i maskopi med honom . 
- Nej , inte alls . 
- Var är han ? 
- Var är han ? 
Varför tog du med dem ? 
Det gjorde jag inte . 
Varför är du här ? 
Vi har inget möte i dag . 
Det här stället har äventyrats , så du måste förflyttas . 
Ni tänkte aldrig skicka mig till Japan , va ? 
Det vet jag inget om . 
Är det farbror Samsiks plan ? 
Nej . 
Du visste ju inte . 
Han skickade hit mig för att det inte är säkert här längre . 
Jag ska förflytta dig . 
Farbror Samsik har förrått mig förut . 
Sineuialliansens uppförandekod Kang Seongmin 
Vem är du ? 
Jag brukade jobba här . 
Vad gör du här ? 
Var är Cha Taemin ? 
Jag letar efter honom . 
Vi hittade de här . 
De har nog tillverkat bomber . 
Jag förstår . 
Gör dig av med dem . 
Ursäkta ? 
Hörde du mig inte ? 
Gör dig av med dem nu . 
Ta en titt på det här . 
- Ska vi bränna det också ? 
Sineuialliansens uppförandekod Kang Seongmin . 
Hallå ? 
Farbror Samsik . 
Det är jag . 
Flyttade du honom ? 
- Det skedde en incident . 
- Vad ? 
Pak Jiwook skickade dit sina män . Och Cha Taemin dödade alla tre . 
Va ? 
Dödade han alla tre ? 
Ja , det gick så fort . 
Cha Taemin misstänker att du försökte döda honom . 
Va ? 
Jag hittade Sineuialliansens uppförandekod , signerad av Kang Seongmin , men Pak Jiwook brände den . 
Signerad av Kang Seongmin ? 
Det hade bevisat att han grundade Sineuialliansen . 
Ja . 
Men han brände den ? 
Ja , framför ögonen på mig . 
Jag är ledsen . 
Okej . 
Bra jobbat . 
Pak Jiwook låter nån skugga oss . 
Liberala partiets ledamot ? 
Ja , han från japanska polisen . 
Vilket mesigt försök att skugga oss . 
Han har även skickat män efter Cha Taemin . Men Taemin ... 
Glöm det . Nu går vi . 
Hur kan koreanskan sjunga så bra jazz ? 
Vem vet ? 
En dag kanske vi slår er i baseboll . 
Den här killen ... 
Du vet Choo Intae ? 
Han som blev skjuten . 
Han har en del anhängare . 
Oroa dig inte för det . 
Det blir inget . 
Jag vet . 
Vi har övat på upploppsbekämpning . 
På amerikanska högkvarteret ? 
Vi genomförde även evakueringsövningar för USA:s ambassad och regeringspersonalen . 
Jäklar . Men det kommer aldrig att hända . 
Men , man ska aldrig säga aldrig . 
Aldrig säga aldrig . Aldrig säga aldrig . 
Krya på dig , herr Choo 
Hur många har dykt upp ? 
Runt 200 . Men folkmassan växer . 
Ilmos sjukhus 
Min far har precis gått bort . 
Partiet måste nu enas för Innovationspartiets framtid . 
Allesammans , det här var ingen olycka ! 
Vi måste ta reda på sanningen ! 
- Ja ! - Ja ! Herr Choo blev mördad ! 
Vi måste ta reda på vem som ligger bakom ! 
- Ja ! - Ja ! Vi måste ta reda på varför det hände ! 
Kom igen , allihop ! 
Vi går till gränden där han blev skjuten ! 
- Ja ! - Ja ! 
Ta tillbaka Choo Intae ! - Ta tillbaka Choo Intae ! - Ta tillbaka Choo Intae ! 
Ta honom tillbaka ! 
Jag åker till sjukhuset . 
Okej . 
Herr Oh . 
Åk och trösta Yeojin . 
Det ska jag . 
Allesammans ! 
Demokratin är död ! 
Ta tillbaka Choo Intae ! 
Av rädsla för att förlora makten dödade de herr Choo ! 
Vi måste gå till botten med det här ! 
Ta tillbaka honom ! Vi måste ta reda på vem som dödade herr Choo ! 
Hur många är samlade ? 
Bekämpar ni upploppet ? 
Det räcker inte på långa vägar . 
Ta tillbaka Choo Intae ! 
- Innovation är vårt hopp ! - Vänta lite . 
- Innovation är vårt hopp ! - Avgå , president Rhee ! 
- Choo Intae som president ! - Choo Intae som president ! 
Ta tillbaka Choo Intae ! - Ta tillbaka Choo Intae ! - Ta tillbaka Choo Intae ! 
Allihop , folket samlas ! 
Vi går ut på gatorna ! 
Kom igen ! 
- Ta tillbaka Choo Intae ! - Förbered eldgivning ! 
- Ta tillbaka Choo Intae ! - Ta tillbaka Choo Intae ! 
Innovation är vårt hopp ! 
- Innovation är vårt hopp ! - Protesten är förbjuden ! 
- Skingra er omedelbart ! 
- Avgå , president Rhee ! 
- Choo Intae som president ! - Choo Intae som president ! 
- Skingra er , annars skjuter vi ! - Ta tillbaka Choo Intae ! 
- Skingra er omedelbart ! 
- Ta tillbaka Choo Intae ! 
Ta tillbaka Choo Intae ! - Ta tillbaka Choo Intae ! - Ta tillbaka Choo Intae ! 
Rhees administration måste avgå ! 
- Avgå ! - Avgå ! 
- Choo Intae ! - Choo Intae ! 
- Lystring , allihop ! 
- Choo Intae ! - Herr Choos dotter är här ! - Choo Intae ! - Choo Intae ! - Choo Intae ! - Choo Intae ! - Choo Intae ! 
Allihop ! 
- Vi måste skingra oss ! 
- Varför ? 
- Nej ! 
- Inte en chans ! 
- Varför då ? 
- Vad pratar du om ? 
Det här är inte vad min far hade velat . 
Det här är inte vad Choo Intae hade velat . 
Han vill inte ha våld ... eller kaos . 
Han stod för vårt folks välstånd samexistens och harmoni . 
Inte ömsesidig förstörelse . 
Min fars död bör hanteras på ett demokratiskt och fredligt sätt . Det är hans önskan . 
Därför måste vi skingra oss omedelbart . 
Det ska inte utövas nåt mer våld . 
- Choo Intae ! - Choo Intae ! - Choo Intae ! - Choo Intae ! 
Ser du ? Inget hände . 
Det vet vi inte än . 
Kang Seongmin vill få igenom lagen om lokalt självstyre . 
Det är din chans att etablera din närvaro . 
Ska jag ska gå emot honom ? 
Du lär dig snabbt . 
Vi vill få igenom lagförslaget så att han kan avancera i Liberala partiet . 
Jag har inget mer att lära dig . 
Genom att motsätta mig framstår jag som en kämpe för demokratin . 
Vi tar en drink till . 
Kl . 21.45 i går avled Choo Intae , Innovationspartiets presidentkandidat . 
Höga popularitetssiffror gjorde herr Choo favorittippad att vinna presidentvalet innan han blev attackerad . 
Det finns misstankar om att Sineuialliansen , en anarkistgrupp , låg bakom attacken . 
Politiska kommentatorer menar att händelsen kan äventyra president Rhees omval . 
Demokraternas kandidat är mycket populär , och många undrar hur händelsen kan påverka presidentvalet . 
Är detta vad jag tror ? 
Ja , de ledamöter som är emot lagändringen om lokalt självstyre . 
Hur många är det totalt ? 
Det är ungefär 20 stycken . 
Så utan deras stöd kan vi inte reformera systemet ? 
Antagligen inte . 
Vad ska vi göra med dessa idioter ? 
Vi kan inte muta dem . 
Tjugo ledamöter är emot lagändringen om lokalt självstyre . 
De utmanar mig officiellt . 
Det är för att vi saknar kampanjbidrag . 
An Yosub försöker ruinera mig . 
Herrn . 
Jag föreslår att du träffar herr An . 
Bageri Sail 
Har du eld ? 
- Jag ? 
- Ja , du . 
Det är jobbigt att förfölja mig . 
Varför kommer du varje dag ? 
- Annars får jag problem . 
- Har du eld ? 
Så du fick sparken på grund av mutor ? 
Ja . 
Här . Det är okej att ta emot mina pengar . 
Gå och ät nåt gott . 
Hur kan du sjunka så lågt och jobba för Pak Jiwook ? 
Återgå till jobbet . 
Ursäkta mig . 
- Jag ? - Han gav dig bröd . 
Farbror Samsik ska träffa Michael Jeong . 
Säg det till din chef . 
Tack . 
Hur mår Yeojin ? 
Har ni pratat ? 
Har du eld ? 
Hur mår du ? 
- Du är tidig . 
- Kom i tid . 
Varför är ni alltid sena ? 
Befälhavaren gav oss sysslor . 
- Vadå ? - Privata ärenden . 
Ta hand om hans växter och keramik . 
Tänk att militärskolan var för det . 
Det är därför vi måste skaka om världen . 
Hanmin . 
Prata inte bara om det . Gör det . 
Va ? 
Prata inte bara om det . 
Varför gör du det inte ? 
Anta att jag gör det . Hjälper du mig ? 
Det beror på vad du gör . 
Vänta och se . Jag ska förändra världen . 
Kom in . 
Herrn . 
Jag får samtal hela tiden . 
Alla gör en stor grej av att be om pengar . 
Kang Seongmin kommer snart och ber om din förlåtelse . 
Vad har hänt med betalningarna ? 
Vet du hur jag framstår om du gör så här ? 
Jag har tänkt göra betalningarna , men ... Jag la dem på is . 
Varför ? 
På grund av den absurda artikeln ? 
Är den absurd ? 
Kan du gå ut ? 
Vad gör du ? 
Jag vet att du misstänker mig . 
Jag erkänner att jag var med i Sineuialliansen . 
Jag formulerade deras uppförandekod . Nej , jag ... Jag etablerade hela organisationen . 
Jag gjorde ett stort misstag som ung . 
Förlåt mig . Men herrn , jag svär ... Jag hade inget med ledamot An Minchuls död att göra . 
Snälla , tro mig . 
Snälla . 
Jag såg Minchul som min egen bror . 
Varför skulle jag döda honom ? 
För att få hans position . 
Nej . 
Jag såg svartsjukan i dina ögon . 
Jag var svartsjuk . 
Svartsjuk på honom . 
Det var jag . 
Så jag såg upp till honom . 
Han uppnådde inte sin dröm . Låt mig förverkliga den . 
Låt mig göra det . 
Snälla . 
Ge mig en andra chans . 
Svär du på att du inte dödade min son ? 
Jag svär . 
Vem dödade då min son och varför ? 
Jag ska ta reda på det . 
Jag ska gå till botten med det . 
Herrn . 
Om Cheongwooförbundet överger mig har jag ingenstans att ta vägen . 
Får jag kalla dig far ? 
Far . 
Jag ska vara lojal . 
Snälla , hjälp mig den här gången . 
Bara den här gången . Skona mig . 
Snälla , skona mig . 
Choi Minkyu lovade att låta dig leda partiet och bli hans efterträdare , eller hur ? 
Ja . Trots det har jag aldrig velat förråda Cheongwooförbundet . 
Hur ska du bevisa det ? 
Jag gör vad som helst . 
- Vad som helst ? 
- Ja , vad som helst ! 
Vill du bli premiärminister ? 
Ta kontroll över Liberala partiet och vinn över 100 medlemmar . 
Sun Wooseok vinner över 40-50 medlemmar i Demokratiska partiet . 
Det finns 20 till 30 oberoende och nyvalda ledamöter som stöds av Cheongwooförbundet . 
Skapa ett nytt parti med de 170 medlemmarna , så kan du bli premiärminister . 
Vad säger du ? 
Kan du vinna över 100 medlemmar ? 
Det kan jag . 
Jag ska få det att hända . 
Oavsett vad . 
Jag ser dig som min son i Minchuls ställe . 
Tack , herrn . 
Kang Seongmin gråter nog vid herr Ans fötter nu . 
Han vet inte att han svalde betet . 
Han är nog tacksam . 
Självklart är han det . 
Han har aldrig drömt om att bli premiärminister . 
Jag har haft honom runt lillfingret sen han var bebis . Vad gör alla amerikanska soldater ? 
Amerikanska soldater ? 
Nåt är på gång . 
Det blev nästan upplopp . 
Ja , men Choo Intaes dotter ... Det räcker . Han har dejtat henne . 
Jag beklagar . 
- Hej . - Hej , Harrison . 
Hörde du ? 
Det är kaos där ute . Vad står på ? 
De yngre officerarna gjorde ett uttalande . 
Om vad ? 
Se själv . 
" Vi motsätter oss splittring , korruption och politik inom militären . 
Alla militärer inblandade i det olagliga valet , samt korrupta generaler , ska straffas . 
Vi kräver en militär reform . Vi kräver bättre behandling av militär personal . 
Vi har vigt vår ungdom till att tjäna vårt land . 
Vår stolthet som soldater har hjälpt oss i svåra tider . 
Vi kräver ansvar av de korrupta generaler som förgör vår stolthet . " 
Du har läst det , va ? Ja . 
Jag skrev det . 
De unga officerarna verkar hålla med om uttalandet . 
Amerikanska arméns högkvarter har ny information . 
Jag håller militären under kontroll . 
Vi kan muta nationalförsamlingen , men inte militären . 
Det såg vi under Japans ockupation . 
Vad för ny information ? 
Militären kan försöka ge förste infaterichefen makten . 
Förste infanterichefen ? 
General Choi Hanrim . Militären litar på honom och han står nära USA:s befälhavare . 
Choi Hanrim ? 
Du träffade väl general Choi på Albrights avskedsceremoni ? 
Ja , det gjorde jag . 
Diskuterade ni statskuppen då ? 
Jag beundrade general Choi mer än nån annan i militären . 
Han hjälpte mig alltid . 
General Choi Hanrim Förste infanterichef 
Han var som en far för mig . 
Minister Kim har så många fäder . 
Det finns många han ser upp till . 
Det är synd att alla hans fäder är döda . 
