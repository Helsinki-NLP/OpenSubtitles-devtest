Jag ska uppdatera dig . 
I morse utsåg drottningen mig till kapten för sin livvakt . 
Låt mig föra dig i säkerhet . 
Hon ska bosätta sig på Broadwater Hall . 
Sofia . Hon ligger bakom allt . 
Besitta varje dödlig sak på ... De ska ta drottningen . 
Hoppas du har turen med dig , Nelly . 
Jag behöver inte tur . Jag har dig . 
Jag tror vi ska stå upp när något är fel . 
Det här är vad vi skickades hit för . Utan för de här stackarnas skull ... Du är min vän . 
Sofia , din far köpte mig ! 
Rasselas är inte mitt riktiga namn . Lord Blancheford gav mig det . 
Mitt riktiga namn är borta . 
Jackson dödade inte min far . Thomas gjorde det . 
- Gjorde han ? 
- Det var han som gav mig idén . 
Jag kan få det att ta slut . 
Isambard Tulley , du ska hängas för dina brott . 
- Stoppa honom ! 
- Jag vet att du är där , Sofia . 
- Ras ! - Du ska inte ... Någonstans . 
Nell Jackson känner till invasionen . 
Vi tar drottningen i morgon . 
Vi ska stoppa dem . 
Lägg undan den , Billy . Du gör mig nervös . 
Hon är sen . 
Det är hon inte . 
Var är vagnen då ? 
Om vi inte tar drottningen här tar Poynton henne . Då invaderas England . 
Då blir det krig och blodspillan , slakt och förödelse . 
Var är hon ? 
Det är snabbaste vägen till Broadwater . 
Hon kommer . Det är bra . 
Har du tänkt på vad du ska säga ? 
Om det blir fel och hon ignorerar dig blir hon kidnappad eller halshuggen . 
Sen invasionen , slutet för England . Världens ... - Du . - Varför inte ? 
Det händer . 
Det är drottningen ! 
Vi rånar drottningen ! 
- Okej . Kör , kör , kör ! 
- Ja . 
- Stå och leverera ! - Leverera ! 
Vi kapitulerar . 
- Va ? 
- Det är skamligt . 
Tänk om hon var en riktig stråtrövare ? 
- Otroligt . Ge mig den . 
- Ja . 
Det är Nell Jackson . Ursäkta att jag kidnappade er , Ers Majestät . Men det pågår en komplott mot er på Broadwater . 
De två drev er rakt in i den . 
Så vi tänkte att det var bäst att fånga dig innan jakobiterna . 
Nelly Jackson ! 
Mr Devereux ! 
Var är drottningen ? 
Jag vet inte . Antagligen i den andra vagnen . 
- Hon använder lockbetesvagnar för att lura folk och för att undvika det här . 
- Vad gör du i den ? 
- Eularia tipsade mig . 
En tom vagn på väg från London är en perfekt flyktväg , för jag är efterlyst nu , tack vare dig . 
Okej . 
Då blir det Broadwater . 
Vi räddar drottningen . 
Hoppas ni har era turbyxor på er . 
Lystring ! Du ... Du är förrädaren ? 
I dag ska du och jag resa till våra jakobitvänner i Skottland . 
Och när Jakob har bestigit tronen kan ditt folk käbbla för din avrättnings skull . 
Arrestera henne . 
Stanna . 
Toppen . 
Sätt fart ! 
Stanna ! 
- Stanna där ni är ! 
- Stanna där ni är ! 
Drottningen är i vårt förvar . 
Våra namn hamnar i historieböckerna . 
Och Poynton ... Du är glad att han hittade dig i London . 
Är du glad att han drog in dig i det här ? 
Ja . 
Så ni är vänner ? 
Har du tänkt om dina fördomar mot honom ? 
Helt och hållet . 
Att skylla omständigheterna på samhället . Yttre influenser . 
Det är en abdikering av vilja . Det gör en till ett verktyg . 
Du låter som ... Fick du den av Poynton ? 
Ta av den . Thomas ... 
Den kan inte tas bort . 
Nej . Sluta ! 
- Vad gör du ? 
- Jag vet inte . 
Jag bara ... Jag måste göra nåt . 
- Jag kände något dåligt . 
Något ont inuti Broadwater . 
Nell bad oss vänta medan hon hämtar Drottningen . 
Det är inte drottningen . Det är nåt annat . 
Jag har en känsla . Jag måste nog lita på den . 
Okej , vi är beväpnade . 
Nell sköter vakterna och jag vet en väg in ... Håll koll på honom , George . 
Kom igen . 
Thomas bär ett hängsmycke . Märkligt lik din ring . 
Det är för att trösta honom . 
Du ville bara ha honom nära när du fick veta att han dödade far . 
År av planering för att nå denna avgörande punkt . 
Drottningen i min makt . England vid mina fingertoppar . 
Allt hänger på de närmaste timmarna . 
Och vi pratar om Thomas ? 
Vagnen till Skottland är redo . 
Den avgår inte förrän du berättar varför Thomas bär ett hängsmycke som inte kan tas av . 
Fadermord vrider och förvrider och märker själen på ett sådant sätt att den kan användas av dem som utövar vårt speciella inflytande . 
Användas ? Istället för att använda energin till att frambesvärja , är det möjligt att helt enkelt dra in den i sig själv . 
I vilket syfte ? När processen är klar blir du omätbart mäktig . 
Permanent . 
Varför har du inte gjort det ? 
Det är något som jag , i mitt nuvarande tillstånd , inte kan göra utan stora risker . 
Men du , med din naturliga styrka och talang , kan göra det . 
Nell Jackson skulle inte betyda något . 
Vad skulle hända Thomas ? 
Han har redan förlorat . Men du kan besegra alla , Sofia . 
Det var du som fick honom att tänka på att döda min far . 
Det hade aldrig slagit honom . 
Du trodde att du kunde leka med oss alla . 
Med mig ! 
Makt , död , förstörelse i min hand . 
Makt , död , förstörelse i min hand . 
Makt , död , förstörelse i min hand . 
Makt , död , förstörelse i min hand . 
Din magi är ingen match för min nu , är jag rädd . 
Man ska aldrig ha något att förlora . 
Det gör en svag . 
Herrn ? Herrn ! 
Två patruller borta . 
- Det måste vara Jackson . 
- Ja . Hörde ni , lady Wilmot ? 
Nell Jackson har bestämt sig för att besöka oss . 
Synd att ni inte får se henne dö . 
Billy , hördu . 
- Ja , vad ? 
- Vi är inte klara . 
- Du har rätt , chefen . 
- Jaså ? 
- Lägg ner vapnet ! 
- Jag trodde du var min chef . 
- Som du håller på . 
- Ja . 
Lägg ner vapnet , sa jag ! 
Undviker konversationen . 
- Har du fått nog ? - Ja , visst . 
Jösses , vilken stor pojke . 
Bäst att Hennes Majestät är tacksam . 
Va ? 
Du är en riktig älva . 
Vi är bra på det här . 
Kom igen då . Är du med mig ? 
Jag är med dig , Nelly . Från början till slut . 
Jag har hört att Broadwater Hall har en fin samling av ... 
- Vad ? 
- Pengar . 
Du klarar dig väl på egen hand ? 
Ja . Jag mår bättre efter skottskadan . Och jag är inte rädd för jakobiter eller vargar . 
- Och efter senaste kidnappningen ... 
Kom då . 
Jag kanske kan hitta nya glasögon åt dig . 
Vad anser du om småstölder ? 
Jag är fäst vid dem . 
Det kommer från honom . Jag känner det . 
Snälla . Inga fler spöken . 
- Han åkallade er för att plåga mig . 
- Vem ? 
Sluta ! 
Tyst ! 
Thomas , det är jag . 
Det är Rasselas . 
Jag ger vad som helst . Sluta hemsöka mig . 
Jag ska berätta hemligheten . 
Jag borde inte ha undanhållit det . Okej . Berätta hemligheten tyst så slutar jag hemsöka dig . 
Amadin . 
Det är Amadin . 
Säg det igen . 
Amadin . 
- Vad är det ? 
- Är det en trollformel ? 
Jag hittade papperen när jag var tio . Det är ditt namn . 
Ditt riktiga namn . Far förbjöd mig att berätta för dig . 
Visste du hela tiden ? 
Jag fick inte berätta ! 
Visste du mitt riktiga namn ? 
Varför ändrade han det ? 
Han gillade det inte . 
- Rasselas . 
- Det är inte mitt namn ! 
- Säg det igen . 
- Amadin ! 
Amadin . 
Han förtjänar det här . 
Det handlar inte bara om honom . 
Vi måste hitta Nell och ta reda på vad som pågår . 
Hon är inte säker . 
Ers Majestät ! 
Jag är Nell och jag är här för att rädda dig . 
Okej . Jag gjorde mig av med alla vakter jag hittade . 
Jag borde kunna smyga ut dig . 
Är du okej ? 
Nell Jackson ? 
Ja . 
Innehållet måste vara värdefullt . 
Tror du ... Jag visste det ! 
Hur fångade du den ? 
- Vad ? 
- Anden inom dig . 
Källan till dina krafter . Hur kontrollerar du den ? 
Det gör jag inte . 
Jag försöker rädda dig . 
Äntligen , Ers Majestät . 
Jag har kämpat genom eld och vatten - för att vara här i nödens stund . - Var är Nelly ? 
Kan du stoppa detta ? 
En strid om kronan ? 
Nationens framtid , världens framtid . 
Tillåt mig , Ers Majestät . 
Isambard Tulley , förmodar jag . 
Du , Nelly Jackson . 
En barägares dotter . 
Tror du att du har nåt att säga till om ? 
Efter allt det där . Fullständigt maktlös . 
Vilken besvikelse . 
Rox , vad gör du ? 
Hängsmycket . 
Du måste vara Poynton . 
Visste du att Thomas dödade din far för att imponera på mig ? 
Det var rätt trivialt , ärligt talat . Men det satte igång nåt . 
Ett gnälligt surr . 
Du , Nell Jackson , är en insekt i ett land av jättar . 
En fluga i tältet hos en general som ska leda sin armé i krig . 
Oviktig . Men jösses , så irriterande . 
Det ska bli ett nöje att slita vingarna av dig innan jag leder en invasion och omformar landet - till det rättmätiga ... 
- Ja . Att göra slut på dig skulle lösa många av mina problem , eller hur ? 
Jag ska ge dig en dålig dag . 
Jag kommer att njuta av att förgöra dig . 
Kan du hålla babblan ? 
Låt oss ta det här utanför . 
Okej . 
Befria mig nu från dolda fiender . 
Oskapa , knyt upp , och lossa banden . 
Möt mig bara , din ynkrygg . 
Tiden kan upphöra och elden fånga natten . 
Försiktigt . Den är ganska stark ... 
Han blir svagare . 
Allt som ligger framför mig att förstöra ! 
Denna dödliga pil , denna säkra förstörelse flyger ! 
Drottningen flyr . 
Skulle inte ni ta över England tillsammans ? 
Kom igen . 
Ers Majestät . 
Överraskning ! 
- Bara lite till . - Thomas ! 
- Roxy ! 
- Nell , det är Thomas . 
Magin kommer från honom . 
Vad är det med honom ? 
Poynton livnär sig på mörkret inom Thomas . 
Formeln kommer att döda honom . 
Din idiot ! 
Kan du inte stoppa formeln ? 
Jag har inget kvar . 
Nell ? 
George ! 
Mr Devereux sa åt oss att gömma oss här i säkerhet . 
Nej , ingen av er får vara här . 
- Det är för sent . 
- Vi går ! 
Nej ! 
Jag tar hand om Poynton medan du får ut drottningen . 
Roxy , snälla . 
Snälla , ta hand om George . 
- Jag kommer att minnas det här , Jackson . 
Jag åker inte utan honom . 
Du kommer att dö . 
Ja , men ... Jag tänkte inte dö i sängen . 
Besvärjelsen stoppar hans hjärta . 
Han behöver hjälp . 
Billy . 
Vi kan inte besegra Poynton . 
Han är för stark . 
Du måste hjälpa Thomas . 
Hur då ? 
Du måste lämna mig och gå in i honom . Bekämpa förtrollningen inifrån . 
Jag har aldrig gjort det . 
Om Thomas dör bryts förtrollningen och Poynton vinner . 
Han får inte dö . 
Men Nelly , du är ju min person . 
Jag vet . 
Vi blir ensamma . Jag vill inte vara ensam . 
Nell Jackson . 
Var är du ? 
Billy ? 
Jag vet inte vad som händer . Tänk om jag inte hittar ut ? 
Vi har inget val , eller hur ? 
Tänk om jag inte klarar mig själv ? 
Det kommer du att göra , Billy Blind . 
Det kommer du att göra . 
Farväl , Nelly Jackson . 
Vänta ! Billy ! 
Nej . 
Mr Devereux ! 
- Mr Devereux ? 
- Fungerade det ? 
Makt , död , förstörelse i min hand . 
Tala med drottningen å mina vägnar . 
Säg att det inte var mitt fel . 
Att vi lurades och tvingades av Poynton , men vände oss mot honom i det avgörande ögonblicket . 
Att det är tack vare oss som ert ingripande lyckades . 
Du fick mig anklagad för mord . Utkastad hemifrån . Min syster likaså . 
Han dödade min pappa . 
Och för att rädda det avskummet förlorade jag precis det viktigaste ... 
" Snälla . " 
Det är väl det du vill höra ? 
Ja . 
Vad sägs om det här ? 
Jag gör dig en tjänst . 
Ja ? 
Jag låter dig gå . 
Låt oss se vad ni två tycker om livet på flykt . 
Det här glömmer jag inte . 
Inte jag heller . 
Billy . 
- Nell ? - Hon är där . 
Nell . 
Vad hände ? 
Nelly ? 
Är det möjligt att bli dubbad till riddare flera gånger ? 
Tja ... Nell Jackson från Tottenham och hennes systrar , Roxanne Trotter , Georgina Trotter , och mr Amadin från Benin . 
Nell Jackson . Jag förklarar er oskyldig till mordet på lord Blancheford och benådar dig och dina vänner från alla brott . 
Sir Charles Devereux . Rikets riddare . 
Du vill visst ha ett citat ? 
Nej , allvarligt , sluta klappa . Tack . 
Nell Jackson . Kliv fram . 
Era ovanliga förmågor har uppenbarligen givits till er för att upprätthålla kronan . 
Vi har hört att ni kan fånga kulor rakt ur luften . Det är dags för en demonstration . 
Vänta . 
- Tre . 
- Nell ! 
Två . 
- Vänta . Förlåt . Vänta . 
- Ett . 
Sluta ! 
Jag är inget billigt trick för sprättar att glo på . 
Du missförstår oss . 
Vi tänker utse dig till kapten för vår livvakt . 
Som den där hemska Poynton var ? 
Det vore en stor ära , som tidigare bara förlänats rikets jämbördiga . 
Det vill jag inte . 
Jag behöver det inte . 
Men tack . 
Du är minsann uppfriskande 
Vad vill du då , Nell Jackson ? 
Har du hört om en pub som heter " Talbot " ? 
