- Där är hon . Isabel ! 
- Jag längtar efter att träffa henne . 
Hon har tur som får dig och David . 
Han blir en så bra pappa . 
Det är inte akut , men jag ser varför hjärtat slår långsammare . 
- Har hon hjärtproblem ? 
Problemet är navelsträngen . Den är virad runt halsen . 
- Herregud . 
- Det kommer att gå bra . 
Gemma är i 39:e veckan och redo . 
- Vi gör ett kejsarsnitt i morgon . 
- Och barnet klarar sig ? 
Jag ska sätta den här monitorn på din mage . 
Är Isabel i nöd skickar den en signal och då tar jag över , annars räcker det i morgon . Gemma ... Det ordnar sig . 
Jag har känt Hana hela livet . Säger hon att det går bra , så gör det det . Jag vet . 
Hon är bäst . 
Du har gjort det så lätt . 
Isabel får en fantastisk mamma . 
Jag tror att hon är livrädd . 
Jag är livrädd . 
Det ordnar sig , Charlotte . 
Du har redan gjort det svåra . 
Du har fått henne att genomgå prenatal vård . Tro mig , de flesta adoptioner går inte till så . 
Jag älskar henne . Gemma , alltså . Det gör jag . 
I morgon överräcker jag Isabel och då har du någon annan att älska . 
Tack . 
Gemma ? 
- Hej . - Jag kommer med gåvor . Kanske landets bästa frukostburritos . 
- De bästa ? - Ja . Och jag borde få dricks . 
- Det här är intressant . 
- Ja , väldigt intressant . De har Tater Tots inuti , vilket jag gillar . Har de ? Jag menade att det var två stycken . Jag är också hungrig . 
Jag tror att du utnyttjar min fångenskap för att umgås med mig . 
- Det är löjligt . 
- Erkänn det bara . 
Jag erkänner att du har lappsjuka och att jag är hungrig . Okej ? Kan du sluta ? Kan jag få en burrito , tack ? 
Okej , vad händer med vårt fall ? 
Ursäkta mig . " Vårt " fall ? 
Ja , bilbomben . Vilka andra fall har vi jobbat med ? 
Det är inte min grej . Mordroteln har tagit över . 
Nej . Jag känner dig . 
Det finns inte en chans att du släpper det . 
Okej , avslöjad . 
Jag bad om rapporten och får en notifikation om den dyker upp . 
Du borde ändå dra nytta av mig . 
Du vet att jag kan lösa det . 
Jag kan göra nytta medan du springer runt och jagar katter . 
Jag skojar , jag vet att du inte gillar katter . - Är det rapporten ? - Nej . - Det är en bröllopsinbjudan . 
- Aj ! Exet går vidare . Inget " aj " . " Ex " är nyckelordet . 
Okej , så du är inte bitter ? Du känner dig inte misslyckad ? Eller dövar smärtan med vem som helst ? Okej . Du är bara glad för deras skull ? 
- Jag är glad för deras skull . - Okej . Jag är så glad för din skull ! 
- Jag gråter inte , du gråter ! - Sluta ! 
Själva ceremonin kommer inte att förändra något . 
Jo , det kommer den ! 
Ceremonier är så viktiga . 
Jag är glad att du säger det , för vi vill att du förrättar vigseln . 
- Det skulle betyda mycket . 
- Ja ! Oj ! Ja . Så klart . 
Ja ! Det vore en ära , ja ! 
- Får jag ta med en gäst då ? - En gäst ? Vem ? Så spännande ! - Jag visste inte att du dejtade . - Jo , och det är en riktig person . Han lever i det här århundradet . Han har bara lite hög profil , och vi är inte redo att gå ut med det än . - Vem ? Kom igen ! 
- När du har tid . 
Du räddades av gonggongen , men samtalet är inte över . 
Navelsträngen är virad runt barnets hals . 
Gemma måste förlösas med kejsarsnitt . 
Om värkarna sätter igång kan det vara för sent . 
Tanken på vad hon ger upp kan ha skrämt henne . Nej . 
Hon fick ett sms precis innan hon försvann . Det verkade störa henne . 
Det har gått två timmar nu . Mobilen går till röstbrevlådan och hon är inte hemma . 
- Hon kanske behöver smälta det . - Inte när barnet är i fara . 
Gemma skulle aldrig riskera Isabels liv . 
Jag förstår . 
Jag har adopterat två barn , det är ett extra lager av oro . 
Det handlar inte bara om barnet . Gemma har blivit en del av familjen . 
- Jag är orolig för hennes skull . 
Jag är också rädd , men för att Gemma har ändrat sig . - Aldrig . 
- Det sa vi första gången också . 
- Det var annorlunda . - Kanske . Jag gillar Gemma , men vi vet hur det slutar . Hon lämnade kontoret . 
Om hon valde att gå , finns det inget vi kan göra . 
Jag hatar att säga det , men han har en poäng . 
Ska vi inte gå ut med en varning ? Jag tycker det . Men vi har en ny chef som " får problem att försvinna " . 
- Så vi får inte orsaka problem ? - Du får inte det . 
Om du efterlyser någon som försvunnit av egen fri vilja , så ... 
Så är jag en känslosam kvinna ? 
- Nej ! Jag värdesätter mitt liv . - Bra . 
Men vill du verkligen reta upp honom ? 
Du har helt rätt . 
" Man fångar fler flugor med honung . " Jag går och häller på honung . 
Espagnol , mi amor ... 
Du ska ju lära dig spanska ! 
Jag var på väg till dig , Batista . - Märkligt . 
- Mustaschen ? Eller hur ? 
Nej , jag var på väg till er . 
Vi kan prata på vägen upp . 
Det är fint utan mustasch . Det ser bra ut . 
- Frun sa att jag rev bebisen . 
- Grattis igen . 
Ni ville träffa mig ? Är det något problem ? Grant har begärt ut en mordakt . Kom förfrågan från MPU eller är din cowboy en cowboy ? 
Jag får återkomma om det . 
Det är Helen . 
Hon gillar musikallåtar . 
Helen ? Ja , jag minns . 
Märklig prick . 
- Jag åker ner igen . 
- Jag följer med . 
Jag ville ha er välsignelse gällande ett fall . 
Vi har en saknad kvinna , gravid , barnet är i fara . 
- Hon är inte efterlyst ? - Nej , inte än . 
Vi försöker klargöra situationen . 
Jag väntade länge på att bli pappa och det gör det än mer värdefullt . 
Som sagt , småbarn kommer först . 
Utfärda en efterlysning . Nu . 
Det finns integritetsproblem , men en adoption kan sluta mycket olyckligt . 
Jag behöver namnet på den biologiska pappan . Jag ordnar en fullmakt . 
Gemma har setts på ett fik i södra Philly . - Så hon gick frivilligt ? 
- Nej . Gemma beställde en ängelshot i kaffet . 
Jag vet , kod för SOS . Hon är i knipa . 
Innan servitrisen kunde skaffa hjälp , tog mannen med sig henne ut . 
- Kameror ? En beskrivning ? - Inga bilder , beskrivningen är vag . 
Barnet överlever inte utan ett kejsarsnitt . 
Samla alla nu . 
Gemma sågs senast kl. 09.15 på en läkarmottagning på Rittenhouse Square . 
- Hon gick inte ut genom ytterdörren . 
- Garaget , då ? 
Hundratals bilar kör in och ut och skyltarna syns inte . 
Många skulle göra allt för ett barn . 
Att ge sig på en kvinnoklinik är vidrigt , men logiskt . 
Mannen måste vara någon hon känner . 
Vad vet vi om henne ? 
Hon är 23 år , född i Pittsburgh . Har inte pratat med sin familj sedan hon hoppade av college . 
Inga sociala medier och inga dejtingappar . 
Bra , men hon hittade pappan någonstans . 
Ja , vi vänt oss till adoptionsbyrån . 
Hans namn finns i papperna . 
- Arbetsstatus ? 
- Hon är säljare på The Punch . De tillverkar kosttillskott till idrottare . 
Vi kollar hennes rundor och stamkunder . 
Vi måste titta på adoptivpappan också - David . Han ville inte att vi skulle leta . Jag är osäker på om han vill ha barn . Han kanske inte vill ha ett barn som inte är hans . 
Vem vill ha ett barn som biologiskt inte är deras ? - Jag menade inte ... - Jag tolkade inte David så . Men vi måste titta på allt . 
Sätt igång . - Jason , mitt kontor . 
Får jag problem för att jag är sarkastisk ? 
Mike tänker som en polis - som ni ska göra . 
Jag jäklas med honom , Nik . Det är allt , okej ? 
Ärligt talat , han stjäl min fru ! 
- Fick du inbjudan ? 
- Ja . Det är bra , Nik . 
Jag är glad för er skull . - Bra . Jag var lite orolig . - För vadå ? Att jag inte har kommit över dig ? 
Jag är lättad . Jag slipper betala underhåll . 
Jag tjänar mer än du , Jay . 
För att du tvingade på mig det här jobbet . 
Ja , ett jobb på MPU , så varför begär du ut en mordakt ? 
Någon utnyttjade oss , och jag vill veta vem . Ja , men det är inte vårt fall . 
Min nya chef friar hellre än fäller . 
Kan du hålla dig innanför linjerna för en gångs skull ? 
Knack , knack . Informationen från adoptionsbyrån har kommit . Den biologiska pappan är en pärla . Vi pratar om snatteri , knarkdomar och han jobbar på ett boxningsgym som Gemma säljer till . 
Han hade ett möte med övervakaren i morse , nära där Gemma togs . 
Messa adressen till gymmet . 
- Stället luktar som en suspensoar . 
- Det är doften av själ . 
Stället har en historia . 
Två Golden Glove-mästare har tränat här . Tredje killen i kön till WBC-titeln i weltervikt . 
- Ser du killen i hörnet ? 
- Är det Avery Hawk ? Ja . Han får Don King att framstå som en mes . 
Är du boxare i Philadelphia äger han dig . 
Jag visste inte att du gillade boxning . 
Jag växte upp med Tyson , Hagler , Hearns , Sugar Ray . 
Kom igen , kolla här . 
Är du redo ? Nej , vänta . Se upp . Ducka . 
- Okej ! Jag tror dig . 
- Kom igen , kom igen . 
Du , Marvin ! Marvin , Marvin ... Var inte asocial . Snälla . 
- Förlåt . Känner jag er ? 
- Philly-polisen . 
Sätt dig . - Jag måste ställa några frågor . - Visst . Fråga på . 
Okej , Gemma Stephenson . 
Varför tittar du på honom ? 
Jag vet att du känner henne . - Visst , jag känner henne ... 
- Mer än så . - Du gjorde henne gravid , Marvin . 
- Saken är den ... - Tog du Gemma för att du ångrat dig ? 
- Nej , nej , nej , nej . 
Vi dejtade , hon blev gravid , hon gjorde ett val . 
Det är lugnt . 
Varför är du rädd , då ? 
Vad gjorde du i morse ? 
Fick du lust att ta ungen tillbaka ? 
Jag svär ! Jag lämnade övervakaren och tog en Uber hit . Jag var sen . Är jag sen får jag sparken och då hamnar jag på kåken igen . 
Men jag kom hit kl. 09.29 och har varit här sedan dess . 
Kan du bevisa det ? 
Hallå , hörni ! Har jag varit här hela dagen ? 
Ja , han har varit här . 
Han spillde kaffe på mina handskar . 
Jag är ledsen för det . 
Igen . - Så vi är tillbaka på ruta ett ? 
- Nej . Det är någon som känner henne och svaret kan finnas i hennes telefon . 
Det tar tid att få ut de uppgifterna . 
Vanligtvis , men jag kanske har en lösning . Bra . Julio Jones ? - Vem ? 
- Din mystiske dejt ? Nej . Varför skulle jag hålla det hemligt ? Jag menar ... 
Okej . 
Min andra gissning - Cory Booker . 
- Ser jag ut att trivas i New Jersey ? 
Är det något på tok ? 
Jag ska gifta mig . 
Varför skulle jag bry mig om vem Jason umgås med ? 
Nikki ! 
Grattis ! 
Spets och bling är inte min grej , men jag älskar bröllop . Jag gråter som ett barn varje gång . Jag vet vad du tänker säga ... 
Att det ser illa ut med en dömd hackare på kontoret ? 
- Hon var min idé . 
Hon är " lösningen " . 
- Toppen . 
Får Gemma värkar innan vi hittar henne kan barnet dö , så ... Jag lovar att inte bryta mot lagen , men jag kanske tänjer lite på den . 
Jag förstår varför ni kommer överens . Tänj , men inte mer . 
Uppfattat , chefen . - Ser du ? Jag är en problemlösare . 
Braun . Om det här tar hus i helvete , får du ta skulden . 
Några framsteg vad gäller barnet ? 
Jag kan följa med ner . Det är tystare där nere . 
- Kan du inte be henne sänka ? 
- Hon jobbar snabbare med musik på . 
Oroa dig inte . Min VPN kommer från Turks - och Caicosöarna . 
Varför därifrån ? 
För om jag inte kan vara där , så kan jag åtminstone vara där . 
Jag vet hur Gemma blev tagen . 
Hon fick ett sms kl. 09.12 . 
" Jag vet att du ljög . 
Möt mig i garaget nu . " 
- Vet du från vem ? 
- En kontantkortstelefon . 
Jag kan inte spåra den . 
När adoptionen inleddes ringde hon Charlotte tre , fyra gånger om dagen . 
För sex veckor sedan dök det här numret upp . 
Det är många samtal . 
Fram och tillbaka . Långa samtal . 
- Du mjölkar ögonblicket . - Det var ett bra ögonblick . 
Okej . Numret tillhörde ... Trumvirvel , tack ? 
Nej . 
- Ett företag ägt av David Ravelle . 
- Charlottes man . - Pågick det något mellan dem ? 
- Ja . Jag grävde djupare . 
Gissa vem som gav Gemma 5 000 dollar varje vecka i sex veckor ? 
Vad betalade David henne för ? 
Gör inte så här mot Charlotte ! 
Jag vet att du inte vill skada henne ! 
Varför har du låst in mig ? 
Gemma kan få värkar när som helst och då kan barnet dö . Ändå vill du inte leta efter henne ? 
Varför har du en engångsmobil ? 
För att skicka ospårbara sms ? Du betalade Gemma för att försvinna , men fick själv ta hand om det . 
Ångrade du dig om barnet eller ville du inte ha det alls ? 
Jag tror att han ville ha barnet . 
Jag har en adopterad dotter . Jag fick panik . Jag fick bara en veckas förberedelser . 
Jag köpte alla böcker och läste dem noga . 
Ja , jag betalade Gemma , men inte för att ge sig av . 
När vår adoption gick i stöpet knäckte det Charlotte . 
Hon ville bara bli mamma . 
Jag betalade Gemma för att stanna . 
Det är olagligt . 
Självklart . 
Vi gjorde allt vi fick göra . Vi betalade alla omkostnader , men jag kunde bara tänka på att om Gemma ändrade sig skulle Charlotte dö . Bokstavligen . 
Så jag sockrade erbjudandet utan att berätta det för Charlotte . 
Jag ville bara att Charlotte skulle vara lycklig . 
Vad är det ? 
Är det Gemma ? 
Det är ett utpressningskrav , de vill ha 100 000 dollar . Du gav någon idén att du skulle betala vad som helst för en nyfödd . 
Vi gör allt vi kan för att hitta Gemma . 
Vi har pratat med hennes jobb , vi kollar alla kontakter . 
Det måste vara någon som kände till adoptionen . 
Släpper de henne om vi betalar lösensumman ? 
Det är alltid en chansning . 
De räknar med att man är villig att göra allt . 
- Jag gör precis vad som helst . 
- Jag vet . Jag säger det här som adoptivmamma , att för det mesta släpps personen fri . Men ni ombeds betala för ett barn som inte är ert . 
Lagen tillåter modern att ändra sig i upp till 30 dagar . 
- Ni kan betala och ingenting få . - Men de släpper Gemma ? 
Kanske . Men det betyder inte att ni får barnet . 
Gemma kommer inte att ändra sig . Hon ligger inte bakom . 
- Det vet du också . 
- Hon säger bara hur det är . 
Vi har sparat och lagt undan pengar till barnet . 
- Vi kan göra det här . 
Vi måste . - Vi kan inte . Jag har spenderat pengarna . Jag betalade Gemma 30 000 dollar . 
- Så att hon skulle göra det . - Hon tänkte göra det ! 
- Hon tog pengarna . 
- Vad skulle hon göra ? 
Hon är ett barn ! 
Trodde du att vi behövde muta henne ? 
Vi gjorde det rätt första gången , och det funkade inte . Jag vet att det är svårt , men vi måste prata om hur ni vill göra när de ger er villkoren för lösensumman . 
Vi hittar pengarna . Det måste vi . 
Jag gör det inte bara för att få Isabel . Jag gör det för Gemma . 
Det hon har gjort räddade mitt liv . Nu måste vi rädda hennes . 
Inspektör Grant . Hollis Braun . 
- Kan vi prata ? 
- Jag är på väg ut . - Kan vi prata på vägen ner ? 
- Hur kan jag hjälpa er ? - Nej , hur kan jag hjälpa dig ? 
Mer specifikt , hur kan jag hjälpa till med Batista ? Hon gör ett bra jobb här . Bara en sak står i hennes väg , och det är du . 
Står jag i hennes väg ? På ditt tidigare jobb tog du genvägar och det belönades . 
- Men här är det ett problem . 
- Handlar det här om akten ? 
Du gör saker som ställer ditt team i dålig dager . 
Nikki är ditt ex . Hon kanske inte känner att hon kan säga det . 
Då gör jag det . 
Du skadar hennes ställning . 
Om det inte förändras , måste vi få det att förändras . 
Ursäkta . Jag bad om en akt , det är allt . 
" Det är allt " ? 
Så det sitter inte en dömd hackare där uppe som gör saker vår avdelning aldrig skulle tillåta ? 
Vi vill alla att Batista ska lyckas , inspektör Grant . 
Försök att hålla dig på din kant . 
Gemmas jobb ger inget . Inga riktiga vänner eller fiender . Jag har gått igenom alla ställen hon levererade till . 
Ingen sticker ut . 
Samma sak med telefonen . Alla blockerade nummer är bara skräppost , indrivare . Det vanliga skräpet . 
- Vänta lite ... - Det låter bra . Betalningarna som David gjorde ... Jag har Gemmas konto här . 
Dagen då hon skrev på adoptionspappren betalade hon 1 000 dollar till Marvin Donald , barnets far . 
- Varför betalar hon honom ? 
- Jag vet inte . Jag kollade inte närmare på honom när han hade alibi . 
- Har du något ? 
- Marvin , din söta lilla lögnare . 
- Jag sa ju att jag har alibi . 
- Även att du var pappan . - Jag är barnets far . - Marvin , lyssna på mig . 
Min chef är på mig , hennes chef är på henne . Jag är inte på humör . 
Det visar sig att när Gemma blev gravid var du i Indiana i en månad . 
Sedan gav hon dig 1 000 dollar . För att köpa en lögn , eller ? Jag kunde inget säga . 
Jag ville träffa mamma och sa till övervakaren att jag hade covid . Det var en lögn , att du var pappan en annan . 
Du bara ljuger . Vill du ha vår hjälp , måste du hjälpa oss . Du måste vara ärlig . Det är enkelt . 
Jag tyckte synd om henne . 
Hon försöker göra det rätta och behövde en signatur för att slippa berätta för den riktige pappan . 
Han skrämde henne . 
Hon sa att han var våldsam . 
- Vem är den våldsamme killen ? - Det sa hon inte . 
Men hon började använda en gymjacka med tigerlogga på . 
Jag tror att det är en av boxarna . 
- Vem är bäst ? - Det är uppenbart . - Creed är bäst . 
- Adonis eller Apollo ? Apollo . Han slog Rocky två gånger . Nej . Första matchen var oavgjord . Det var uppgjort . 
Rocky vann båda matcherna . 
- Jag håller inte med . Vem gillar du ? 
- Adonis . Han studerade sin far , Rocky tränade honom . 
I vilken värld slår Michael B. Jordan Carl Weathers ? 
Kolla på " Rocky " ! 
Det är min åsikt . 
- Va ? Jag pratar ! 
- Här är listan . Alla som har köpt en jacka , men den kom inte från mig . En sak ? Smyg dig inte på folk så där . 
Gå nu . 
Du har gjort tillräckligt . Ska vi ta alla på listan , en efter en ? Jo , vi har ju hela dagen på oss . 
- Du får inte ringa i klockan ! - Kan jag få er uppmärksamhet ? 
Vi är från polisen . 
En av er snygga , unga boxare gjorde tillskottsflickan gravid . Vem ? - Griper ni folk som har sex ? - Nej , men du är rolig . Du borde prova ståuppkomik , för din boxning suger . Någon måste erkänna , annars blir det inte mer träning i dag . 
Eftersom fyra av er ska tävla i kväll , så suger ju det . Jag skickar runt ett foto . En av er måste erkänna . 
Som han sa , sex är inget brott . 
Det är sex . 
Det är inte olagligt . Vi vill bara veta vem . 
- Namn ? - Dante D ' Andrea . 
- Ja , han är med på listan . - Berätta om dig och Gemma . 
Heter hon så ? Jag har sett henne , men känner henne inte . 
Hoppas att du är bättre på att boxas än att ljuga . 
Jag tror att det är han . Gemma sa att han var en mobbare , en osäker kille som vill verka tuff . 
Hon sa att hon aldrig hade gillat honom . 
Sexet var hemskt . Slöseri med tid . 
Våld mot tjänsteman . Ger det två år ? 
Nej , upp till 40 år . Jag kan hjälpa dig , men du måste hjälpa mig . 
Du måste börja prata . Okej ? Jag dejtade Gemma , men visste inte att hon var gravid . 
Sedan såg jag efterlysningen och räknade efter . Jag sa inget , för jag visste vad ni skulle tro . 
Jag ska säga vad jag tror . Du sms:ade henne i morse . 
Vi såg sms:et . Okej ? 
Hon ljög om något , eller hur ? Du bad henne träffa dig och sedan tog du henne . 
- Du vill ha snabba pengar , eller hur ? 
Jag har vunnit tre matcher . Vinner jag i kväll blir jag tät . Mitt sista erbjudande : 
Tala om var Gemma är just nu så får du boxas när du kommer ut igen . Hur ska du ha det , Dante ? 
Vill ni veta om jag är pappan ? Ja , troligen . 
Men jag har inte sms:at och att göra någon gravid är inte olagligt . 
Jag är ledsen att jag slog dig , men det är inte mig ni söker . Okej . Okej . 
Vi hade inget på honom , men fick söka igenom hans ställe . 
- Det gav inget . 
- Vi vet att Gemma inte är där . 
Du är arg för att du fick en smäll . Det är inte mitt fel att dina reflexer är långsamma . 
Tror du Nikki vet att hennes nästa äktenskap blir sämre ? 
- Rent atletiskt , alltså . - Är du färdig nu ? - Hej , Nik . 
- Vad har hänt ? 
- Inget . 
En olycka . - Han glömde ducka ! 
- Hittade ni barnets far ? 
- Han heter Dante D ' Andrea . 
Vi hittade inget hos honom . Säg att ni hade skäl att gå in i hans bostad . 
Han slog Mike i ansiktet ! Vilket är ... ett skäl . 
- Och han är nog den skyldige . 
- Vi börjar få ont om tid . 
Jag vet . Överlämnandet sker på matchen i kväll . 
- Charlotte gör det . 
- Och då tar vi honom . 
Det är bäst , för enligt monitorn blir hjärtfrekvensen svagare . 
Om vi inte hittar Gemma i kväll kan det vara för sent . 
- Försöker du gömma dig för mig ? - Nej , det vet jag att jag inte kan . 
Helt rätt . 
Vad gör du ens här ? 
Du går inte upp i ringen i kväll . 
Det här är mitt event och du ska veta att det är över för dig i Philly . 
- Jag vet att jag klantade mig . - Som om det var en olycka ? 
Du behövde bara förlora , men slog min kille medvetslös . 
Vet du hur mycket jag satsat på Kwan ? Det var dumt gjort . 
Du visste att jag satsade på den andre . Jag har en plan . Du ska få tillbaka allt i kväll . 
- Du tjänar inte 100 000 på matchen . - Nej , du får dem innan matchen . Jag vill bara att du behåller mig på kortet . 
Dödar du mig nu får du ingenting ! 
Jag har en plan . 
Hawk låter mig vara om jag betalar honom . 
Han får sina pengar och jag drar härifrån . 
Jag bryr mig om dig , Gem , men jag hade inget val . 
Jo , det hade du ! 
Jag sa nej ! De är bra människor . 
- Jag behöver bara ett par timmar . 
- Vattnet har gått , Dante ! 
Barnet är på väg , och om jag inte får vård nu kommer hon att dö . 
Det vill du inte . 
Hon är din ! Jag ringer 112 så fort det är klart . Bara ... Om jag släpper dig nu dör jag , så snälla , håll ut lite till . 
Vi måste veta vem vi har att göra med . 
Jag hittade Dantes senaste match . 
Någon hade lagt upp den här . 
Motståndaren var Kwan Ju-Won . 
Det skulle vara en enkel match för Kwan , men se vad som händer . 
- Jag förstår Gemmas rädsla . - Kwan ligger fortfarande i koma . 
Meddela alla att de ska närma sig med försiktighet . 
- Jag har ritningarna över arenan . 
- Okej . Vi går igenom planen . 
Så fort första matchen börjar lägger Charlotte pengarna i en väska och går in på arenan . 
Inga poliser syns till . 
Mike och Jason är i säkerhetsrummet . 
Vi har ögonen på pengarna , på Dante , på allt . 
Charlotte lägger pengarna i ett brandskåp och går därifrån . 
Vi har uniformer på plats och vi har vårt hemliga vapen . 
Kidnapparen tar pengarna , men vi tar honom inte förrän han leder oss till Gemma , för vi spårar väskan . 
- Han drar nytta av folkmassan . 
- Vi följer pengarna . 
Han har rocken på och är tejpad . 
Vänta , vänta . 
Kolla hur rocken sitter på honom . - Han är en lättviktare . 
- Väger han för mycket ? Jag tror att vi har blivit lurade . 
Vad gör du ? 
Enligt Kemi är pengarna kvar . Han tejpade inte händerna , han tejpade fast pengarna på kroppen . 
Den misstänkte är Dante D ' Andrea . Han måste hållas under uppsikt . 
Han tog pengarna från andra sidan . 
- Vad finns på andra sidan väggen ? 
- En servicekorridor . En väg leder till östra trapphuset , den andra till nedre hallen . 
Nedre hallen . Vi delar på oss . 
Dante tänkte aldrig boxas . 
Det var en skenmanöver . 
- Ta upp säkerhetskameran igen . 
- Charlotte ! 
Där ! Alla enheter , en civilperson är på väg mot servicekorridoren . Vit kvinna , 35-40 år , med rutig scarf . - Han är i den nedre hallen . 
- Jag är på väg . Vänta ! 
Han såg poliserna vid nordvästra utgången . 
Han går tillbaka mot Mike . 
Jag ser honom inte . Polis ! Dante , stanna ! 
- Han springer österut . 
Jag kommer från andra sidan . 
Han är i förrådet i östra korridoren . 
- Hallå ! Dante , hördu ! 
- Låt mig gå härifrån . 
- Rör dig inte . - Var är hon ? 
Lyssna på mig . Släpp henne , så pratar vi . 
Dante , vi kan hjälpa dig . Det är kvinnan som ska ta hand om ditt barn . - Hon förtjänar inte att bli skadad . 
- Håll käften ! Jag går härifrån nu . - Okej , okej . 
- Lägg ner vapnen ! 
Lägg ner dem ! Sparka bort dem ! 
Ser du ? Jag ska inte skada dig . 
- Ta det lugnt . - Jag ville inte det här . 
Jag svär . Jag ska släppa dig . Så fort jag kommer till dörren . 
- Är du oskadd ? - Ja . Hallå ! Dante ! Håll dig vaken . 
- Få hit en sjukvårdare nu ! 
Vi får inte något ur honom . 
Han är den enda som vet var Gemma är . 
- Herregud ! 
- Vad är det ? 
Den larmade . 
Det är dags att föda . 
- Vi har hittat hans bil . 
- Var har han henne ? 
- Vi ser inget här . - Det ni inte kan se då ? 
- Kan du utveckla det ? - Ge mig VIN-koden . 
Har du den ? Då så . 
- VIN-koden kommer här . 
- Ge mig den , tack . - Ja , självklart . 
Bilar är numera som mobiler på hjul . 
Datan laddas upp automatiskt upp till platser du inte vill känna till . 
- Så du får platsdatan ? 
- Då måste jag hacka OnStar . Men här är alla platser där bilen har stått sedan Gemma togs . Parkeringskameran sparar datan . Det är Barella ' s , den kan du ta bort . Förlossningsläkarens kontor , inte det . 
Okej , och det är fiket som kommer härnäst ? Jag vet inte var det är . Bilen återvände hit efter samtalet med Dante . - Kan du få fram en adress ? 
- Nu ber du om mirakel . 
Jag utför mirakel . 
Skicka bilden till mig . - Härligt . - Vi tar fram bilden . 
Jag ska förstora det där . 
Titta på skylten i bakgrunden . 
Är det koreanska ? Hur hjälper det ? 
Kwan , boxaren som Dante försatte i koma , bor i Koreatown . Dante visste att hans lägenhet stod tom. 
- Ge mig hans adress ! 
Bra jobbat ! 
- Snyggt . 
Bra ställe att hålla gisslan på . 
Okej , se upp . 
Ur vägen . 
- Vad gör du ? 
- Skjuter av gångjärnet . 
Med en gravid kvinna och eventuellt en bebis där inne ? 
Stolt ? Mitt sätt hade också fungerat . 
Sätt fart nu ! 
Gemma , Gemma ... Allt kommer att bli bra . 
Barnet ! 
Nikki , vi är inne . Det händer definitivt nu . 
Läkaren är på väg . Titta på mig . 
Allt kommer att bli bra . 
- Ge mig lite utrymme . - Jag är här , Gemma . 
Förlåt ! 
Jag är så ledsen ! 
Vi hinner inte ringa efter ambulans . 
Kom in . 
Tack , Hana . 
- Hon fick bort navelsträngen i tid . 
- Vill ni hålla er dotter ? 
Tack , Gemma . 
- Här . 
- Tack . 
Du måste ha älskat att se henne hålla barnet i dag . 
- Ja , det var otroligt . - Var det det ? 
Jag minns första gången jag höll Sidney . 
Vi tog hem henne och hon var så rädd . 
Jag höll henne i mina armar . 
Det lugnade henne , men det förändrade mig . Det förändrade allt . 
Nu är Keith borta och Sid iväg på sitt håll . 
- Jag saknar det . 
- Jag vet . 
Det är okej . Det är så cykeln ser ut , men jag saknar det . 
Det är grejen med cykler . Det finns alltid en chans att påbörja nya . Det var aldrig något vi bestämde oss för . Det var kaos med Keith , och det räckte men vi kanske borde överväga det . 
Ska vi ta in på den vägen ? Påbörja vår egen cykel ? 
Jag vet inte . 
Vi kanske kan börja med bröllopet och ta det därifrån ? 
Okej . 
- Okej . 
Är det fel att vilja att någon annan blir tagen i morgon ? - Ja , det är väldigt fel . 
- Ja . Men jag hade kul i dag . 
Det var en sjujäkla dejt . 
Näta gång du vill träffa mig , så kan du bara fråga . - Jag gillar inte bondage . - Sätt dig . Bossig ! 
- Tack . 
- Du behöver inte sätta fast den . 
Du var inte så besvärlig i Kandahar . 
Du var gift och jag uppförde mig . 
Just det , ja . 
Jag borde gå . 
Jag måste gå nu . 
Den där bilbomben , då ? 
Du hade rätt , jag lider av lappsjuka . Okej , så här är det . 
Vår nye chef är besvärlig . 
Han var arg för att du var där . 
Nikki bad mig backa , så jag backar . 
- Hon ska gifta sig med en annan . 
- Vad fan ska det betyda ? 
Den Jason jag kände skulle aldrig låta en chef stå i vägen . 
- Okej , du vinner . 
Varsågod . 
- Tack . - Du behöver ett användarnamn och ... 
- Jag är redan inne . 
Jag tillbringade hela dagen på MPU . 
Det är en vanesak . Ärendenummer ? 
Ja , det är Hotel-Oscar Monster-26984 . 
Vad är det ? 
Det utlöstes ett virus när jag öppnade filen . 
Filen är vitlistad . 
Någon vill verkligen inte att du ska se filen . 
En utöver Nikki har sagt åt mig att backa . 
Det är överintendenten . 
Vad vill Hollis Braun att jag inte ska se ? 
