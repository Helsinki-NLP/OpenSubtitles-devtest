TIDIGARE I SERIEN ... 
Bob blev nog glad när han hörde vilken loser jag visade mig vara . 
Att ha fått sparken gör ingen till loser , Tony . 
Att därför sura och överge familjen , gör det . 
- Du kan begå ett misstag ! 
- Så som du ! 
Tilly föddes mindre än nio månader efter att ni gifte er . Jag vet vad det betyder . 
Vi hittade Van . Han är på ett flyktingläger i Malaysia . 
Jag känner en malaysisk man . Han kanske kan hjälpa er , men han tar betalt . 
- Poppy , titta , han hämtade din byst . 
- Vad ska du med den ? Det brinner ! 
Vår Stirling brinner ! 
- Vad är ditt problem ? 
- Du borde inte ha kysst honom . 
De har inte vad du har , men de verkar trevliga . 
Vi kan göra det bättre . 
Kvinnor åker inte till rymden längre . 
Bättre att bli skönhetsdrottning , va ? 
- Ge den tillbaka ! - Vill du ha den ? 
- Kom och ta den . 
- Ge min bräda tillbaka ! 
- Vad gör du ? 
- Vad gör du ? 
- Du kan inte ens köra . 
- Du ska få se . 
- Du skulle bara våga ! Hallå ! 
- Stanna ! 
Du kör för fort . 
- Jag försöker ! 
- Hårdare ! 
Nej ! 
Är du okej ? 
Backa . 
Bakåt . 
Chook dödar oss . 
SCARBOROUGH BEACH SJUKHUS 
Det här är skit . 
Era barn stal bilen . 
Det är en brottslig handling . 
De kan hamna i belastningsregistret . 
Kom igen , Rocco . 
Det var ett misstag . De är bra ungar . Du känner dem . 
Jude , bra ungar stjäl inte bilar . 
Du är pappa . 
Kan du inte ... Jag skulle älska det om du kunde få det att försvinna . 
Jag skulle älska att hjälpa dig . 
Okej . 
Jag skulle älska att inte måsta åka hemifrån om kvällen för att föräldrar inte har koll på sina barn . 
- Rocco , jag ... - Va ? 
Att sändas ut till en olycksplats och inte veta om jag får sopa upp döda kroppar . 
Om bilen hade träffat trädet lite annorlunda , skulle du behöva en begravningsentreprenör . 
Men ja . Visst , Tony . 
Jag ska få det att ... försvinna . 
Det kommer aldrig att hända igen , Rocco . 
Du , han har ju rätt . 
Jag minns inte att vi tvingat henne ut i natten för att bete sig som en idiot . 
Det som hände borde inte ha hänt . 
Vi har varit distraherade . 
Är du nöjd , va ? 
Det är inte jag ! 
Min bräda ! 
Varför har de gjort så ? 
- För att hålla henne borta från stranden . 
- Åh , Mia ! Älskling ! 
Mia . 
Såg du dem inte ? Eller hörde dem ? 
Ringde du polisen ? 
" Är du okej , Tilly ? 
Hoppas du inte oroade dig , Tilly . " 
Jag är okej , mamma . 
Tack , pappa . 
Jag vet att ni tänker på mig . 
Han behöver grön olja . Det läker fortare . 
Här , jag har . 
Tack . 
- Nej , jag är okej ... 
- Bråka inte . 
Det blir varmt idag . 
Ni kommer att ha fullt upp . 
Har du ringt ? 
Jag pratade med den malaysiske mannen . 
Är han från ambassaden ? 
Är han här eller i Malaysia ? 
Det enda viktiga är pengar . 
Fem tusen säger han . Jag garanterar att er son kommer ut ur landet . 
Därefter blir det en ny betalning . 
De vet inte ännu hur mycket . 
Ja , jag ska göra en kassett till dig . Alla hitlåtar . 
" Macho Man " , " YMCA " . Okej ! 
Det vore fint . 
Vad har du råkat ut för ? 
Pappa ? 
Pappa ! Vad gör du ? 
Vad gör den där på min gata ? 
Jag hörde om mitt barnbarns olycka - från matvagnen ! 
- Det är olagligt att parkera här . 
Du har tur att min man inte är hemma ! 
Jag går till fullmäktige . 
Jösses , Bob ! Du välte soptunnorna . 
Någon måste ta kontroll över familjen - så nu flyttar jag in . 
- Kan jag få betalt ? 
Jag går efter nycklarna och kör dig till stranden . 
- Nej ... 
- Pappa ! 
- Jag går ingenstans . 
- Vad gör du ? 
Du måste ta huvudet ur arslet och skaffa dig ett jobb - så att min dotter kan vara en god mamma . 
- Åh , visst . 
Men när jag hade ett jobb gillade du inte det heller , va ? 
- Avgiften är fem dollar . 
- Nej , det var ditt agiterande . 
- Ja , ditt agiterande . - Mitt agiterande ! 
- Det ogillade jag . - Jaha ... 
Fackföreningslarvet . När du borde ha varit hemma med dina barn . 
- Vad vet du om det ? 
- Gå inte ifrån mig . 
Hon är vuxen och gör som hon vill , Bob . 
- Hallå ... - Betala honom . 
Hallå , lyssna ! 
- Jag vill träffa Mia . 
Hon behöver mig ... 
- Hon behöver vila . 
Kom inte in i mitt hus . 
Du får göra om den . 
- Vad ? 
- Stirling . 
Karlen som du grillade på gårdagens fest . 
Mamma skulle vara stolt . 
Du är inte här för ett politiskt uttalande . - Du är här för att få en utbildning . 
- Jag är inte den som behöver utbildas . 
Jag ska säga dig en sak . 
Den smartaste mannen jag känt dog i fängelse . 
Han fattade inte , att göra vita arga får dem inte att lyssna . 
Hej . Ja , din son är här . 
Ja , han har stora planer för veckoslutet . 
Den där bysten du gjorde . Kan du lära mig att göra en ny ? 
Ja ! 
- Ja ? 
- Ja . 
Men ... din pappa och mamma ? Är de hemma ? 
Nej . 
Lördagar fixar hon håret . 
Stort projekt . 
Vad han gör vill jag inte ens veta . 
Eller jag vet , men jag önskar att jag inte gjorde det . 
- Du först . 
- Okej . 
- Får jag ? 
- Okej . 
Tack ! 
Försiktigt . 
Ta-da ! Finrummet . 
Vi gör det här . 
Ja . 
Nej , jag förstår . 
- Vad bränner vid ? 
- Han är redaktören . 
Jag vet inte om det är rätt tillvägagångssätt , Wayne . 
Om du ger mig numret , kan jag ringa till honom . 
Okej . Tack . 
Jag försökte slipa bort det som de skrev på brädan . Det sitter för djupt . 
Någon dog på sjukhuset på grund av strömavbrottet . 
Tänk om det hade varit Mia . 
Wayne vill att jag håller det ifrån tidningarna . 
Det förstår jag . 
Han säger att sjukhuset också vill undanhålla det . 
Han måste förstå - att det får konsekvenser ... - Om strejken hade lösts , 
- skulle vi inte ... - Så det är mitt fel , va ? 
Tony , det menar jag inte . 
Det här är inte mina mäns fel . 
Om företaget behandlade oss rättvist , 
- skulle vi inte ... - De är inte dina män . 
Älskling , det är inte din kamp . 
Mia ? 
Kom igen ! 
Vågorna väntar inte ! 
Jag är trött på Stirling . 
Vad är så speciellt med honom ? 
Han seglade bara nedför en flod . 
Har du hört om slaget i Pinjarra ? Nej . 
Stirling vann det . 1834 , 25 män . 
De steg upp två timmar före gryningen för att fienden inte skulle se dem komma . 
De smög ner längs Murray . 
Stirling var ledaren , men han gick knappast först . 
Ja , vi pratade om det i skolan . 
Var det inte någon som dog ? 
Jo , en polis . 
Och cirka 80 Pinjarrabor . 
Också kvinnor och barn . 
Varför gör vi då den här bysten ? 
Det gör vi inte . 
En mellanöl , tack . 
Tony tamejfan Bissett . 
George . 
Jag saknade dig på mötet . 
På alla 17 möten , faktiskt . 
Jag gillar inte möten . 
Ja , du missade inte mycket . 
Bara skalliga karlar och ölmagar . 
Hur i världen ser du fortfarande så bra ut ? 
Är du okej ? 
Jag är sjuk på grund av öknen . 
Vi kan inte prata om det . 
- Vi skrev på det där pappret . 
- Jag bryr mig inte . 
De brydde sig inte om oss när de utsatte oss för radioaktivt nedfall med de där testerna . 
Jag pratar med en jurist . 
Men vi behöver siffror om vi ska sätta dit dem . 
Det är brittiska regeringen , 
- för Guds ... - Du , lyssna på mig . 
Vad du än gör , vill jag inte vara inblandad . 
Jag har aldrig pratat om det , och tänker inte börja nu . 
Du klarar det , miss Universum . 
Miss Sovjetunionen är förstasidesstoff och allt populärare på grund av entusiasmen för allt som är australiskt . 
Katrina Munro , Kanal Två , Perth . 
Okej , damer , vi gör en rad . 
Ge mig kapporna . 
Skynda på . 
Tack . 
Tack . 
- Jag ger henne en åtta . 
- Såja . 
Nio . 
Hon tappar poäng för heldräkten och håret . 
Jag föredrar blondiner . 
Vem bryr sig . 
Jag säger inte nej till någon av dem . 
Ställ miss Sovjetunionen i mitten . Jag gör det värt din möda . 
Ursäkta , ett ögonblick , herrar . 
Vänta lite ! 
Fort . 
Flytta på er ! 
Vinka och säg , " Hej Perth ! " 
Hej , Perth ! 
Att filma festen var mycket smart . 
Hon är en vanlig tjej . 
Hon äter deras mat , leker med deras barn . 
Nu när hon är på toppen måste hon hållas där . 
Visa lite personlighet ! 
Har du varit i militären ? 
Vietnam . 
Jag lärde mig hålla ciggen så här på grund av regnet . 
Nu är det främst en vana . 
Min son är i armén i Afghanistan . 
Han är ingenjör , men snart blir det krig . 
Det är alltid krig . 
Tack , herrar . 
Har ni frågor till flickorna ? Nu har ni er chans . 
Bra . 
I morgon kväll får jag ta med en gäst . 
Jag känner mig som Askungen . 
Guvernörens bal . 
Bara rika människor . 
Ingen vanlig kostym . Smoking . 
Dansar du ? 
Som Nurejev ? 
Ungefär . 
Vad ? 
Gäller ditt erbjudande ännu ? 
Ja . 
Jag har ett jobb , bara så du vet . 
Vill du ha en medalj ? 
Mia ? 
Mia är i duschen . 
Hon är där i en evighet , så ... 
Är hon okej ? 
Mia är alltid okej . 
Om hon inte pratar med mamma , kommer hon inte att prata med dig heller . 
Kanske du borde försöka . 
Varför skulle jag försöka få Mia att känna sig bättre ? 
Kanske för att hon är din syster . 
Och inget illa har hänt dig . 
Tror du verkligen det ? 
Jag trodde att jag höll på att bli sjuk , och ville inte smitta din mamma . 
- Var är Mia ? 
- Var tror du ? 
Vad är det med dig ? 
Du låter åtminstone frisk . 
Har det blivit bättre ? 
Han har sovit på soffan . 
Han gick ut i går . 
Vem vet vad han gjorde , eller var . 
Jag menade Mia . 
Åh , naturligtvis . 
Hon äter inte . Hon pratar inte . 
Hon kommer inte ur sängen . 
Alla flickor går djupt . 
De är som valar , de dyker ner . Man ser dem inte på flera dagar . 
Pojkar hoppar runt dig som idiotiska delfiner . 
Jag är portad från Chez Bissett . 
- Den vanliga ? 
- Härligt . 
- Hur har du haft det ? 
- Bra . Jäktigt . 
- Jag bjuder . 
- Åh , nej . 
- Tack ! 
- Och den här . 
Jösses . 
Våra besparingar . 
Fem tusen för Van . 
Sandy ... 
Tack vare dig kommer vi att vara tillsammans . 
Man kan inte köpa sig in . 
Eller man kan , men en biljett kostar tusen dollar . 
Det är sådant folk där i kväll . 
Köper du dig en bättre danspartner ? 
Alla som är någon kommer att vara där . 
Murray Doull är där . 
Får jag fem minuter med honom , får jag honom att investera . 
Vad hade du gjort om jag inte var här ? 
Du är alltid här . 
Kul att du märkt det . 
Tänker du inte säga något ? 
Var försiktig . 
Jag tror Murray gillar lustjakter mer . 
Eller är det världens vackraste kvinna som du oroar dig för ? 
Jag oroar mig för dig . 
Jag klarade mig ut ur fårklippningen och armén oskadad , - Ja , för att du ville ut , inte in . 
Alla vill inte stå utanför och röka gräs och dela på grönsaker . 
- Dessa människor ... 
- De har pengar att ta mig till nästa nivå . 
Nästa år är jag på gästlistan . Inte bara någon annans gäst . 
Efter i kväll är allt annorlunda . 
Titta inte upp . 
Folk med makt tittar bara på sin nivå . 
Eller ner på vad de vill ha . 
Du måste veta din plats . 
Spela din roll . 
Det är teater . 
Du behöver bara spela teater . 
Vem vill du att jag ska vara ? 
Vad gör du här ? 
Pressen har inte tillträde . 
Han är med mig . 
Du måste mingla . 
Bra idé . 
Nu ska vi träffa stans mest inflytelserika man . 
Mick Bissett . 
Murray Doull . 
Jag tänkte att ni herrar vill träffa blivande miss Universum . 
Godkväll . 
Miss Sovjetunionen , naturligtvis . 
Frank har sett till att alla vet dig . 
När Frank snappade upp historien , hade den redan varit i medierna runt om i världen . 
Frank måste förstå att nyheterna förändras . 
Sovjetunionen är på gränsen att invadera Afghanistan , men en skönhetsdrottning på grillfest är det som intresserar tittarna . 
Vad gör dig till expert i frågan ? 
Svetlana är min historia . 
Hon är min skapelse . 
För två dagar sedan var hon ingen . Nu är hon favoriten . 
Och tävlingen har inte ens börjat . 
Mitt företag , Bissett Star Broadcasting , kommer att revolutionera mediabranschen . 
Nu dansar vi . 
Du har rätt . 
Man kan inte gå på hårt nog med så rika män . 
Man måste spela svårfångad . 
Tror du att jag är din skapelse ? 
Att jag inte vore något utan dig ? 
Du måste erkänna att för några dagar sedan var du ingen . 
Och nu ... Alla tittar på oss . 
Tittar de på oss ? 
Se dig omkring . 
GUVERNÖRSPALATSET VÄLKOMNAR MISS UNIVERSUM 
Du har fel . 
Det är hon som har makten . 
Du kunde ha varnat mig . 
Det är roligare så här . 
Potatis till alla ! 
Ha en trevlig kväll , pojkar . 
Jag tar pengarna också . 
Lam , nej . 
Ni kan väl gå på bio , va ? 
Jag bjuder . 
Jag vill inte gå på bio . 
Jag vill ha en ny bil . 
Är det allt ? 
Jag kommer tillbaka en annan gång . 
Binh , nej ! 
Hallå , ge dem tillbaka . 
Ska du slåss med oss alla ? - Binh ! - Va ? 
- Kom igen ! - Kom . 
Ja , göm dig bakom mamma . Fegis ! 
- Nej , Binh ! 
- Kom igen ! 
- Hallå ! Hallå ! - Lam ! 
Kom hit ! 
Slåss inte . 
Gå ! 
... loser ! 
Vi stänger tidigt ! 
Vi går till templet imorgon . 
Min son , vad tänkte du på ? 
Vi går hem . 
Bra ! Snyggt kast ! 
Mia vill inte ha den , så någon borde äta den . 
Hon måste ha det bra om hon säger nej till shepherd ́s pie . 
Barn ! Läggdags . 
Barn ! 
Som barn ville jag bara ha en normal familj . 
Nu vill jag att mina barn har allt som jag aldrig hade . 
Sedan händer allt detta , jag får det här jobbet och jag tror ... Jag tror jag är bra på det . 
Jag har inget emot långa dagar eller bollande . Jag ... Jag oroar mig att jag inte finns där för dem . 
Jag jobbade , och du blev ju okej . 
Det blir dina barn också . 
Jag vet inte vad jag ska göra med Mia . 
Frågar du mig ? 
Vad skulle du göra annorlunda ? 
Inget , du är perfekt . 
- På allvar , pappa . 
- Jag menar allvar . 
Jag tycker du är lysande . 
Fråga inte vad jag skulle ha gjort annorlunda . 
Det måste ha varit svårt att växa upp utan mamma . 
Åh , jösses . Jag vet att jag inte var perfekt . 
Kanske jag kom hem sent , men du visste att jag skulle komma . 
Varje kväll var jag hemma . 
Det är du också . 
Var är din skugga ? 
Han letar efter bilen som förföljde oss hit . 
Blev vi förföljda av en bil ? 
Det finns alltid en bil . 
Du dansar bra . 
Finns det inte många som dansar bra där hemma ? 
Jag vet hur det är . 
Det fanns inte många där jag växte upp . 
Här i stan finns det fler . 
Här finns mer av allt . 
Hallå ? 
Hallå ? 
- Jag lägger på . 
- Det är jag , Niki Lauda . 
Mia , du kunde ha dött . 
- Du kunde ha dödat oss båda . 
- Men jag gjorde det inte . 
Jag är ledsen för krocken och kyssen ... 
Jag är så ledsen för alltihop . 
Mia ? 
Mia ? 
Mia , sluta lägga beslag på badrummet . 
Andra behöver också använda det . 
Mia ... 
Pappa ! 
Vad är det som händer ? 
Hon behöver sin mamma . 
Det är bra nu . 
Allt kommer att bli bra . 
Vill du prata om något ? 
Var jag ett misstag ? 
Låt mig berätta en historia . 
Jag träffade din mamma när hon började jobba på fabriken . 
Jag var lärling och hon hade ett jobb på kontoret . 
Jag hade just fått mitt körkort och ville bjuda ut henne i bilen jag köpt för alla mina besparingar . 
Men din morfar lät inte henne åka i bilar med pojkar . 
Särskilt inte med en fackföreningsfantast . 
När vi började träffas måste vi ta bussen . 
Tidtabellerna var hemska . 
Det gick en buss till biografen varannan timme på veckosluten . 
Det jag försöker säga , älskling ... är att ingen väntar i två timmar på en buss ... av misstag . 
Enligt NASA har Skylab , den för tillfället obemannade rymdstationen hamnat i en sjunkande omloppsbana . 
Detta är det senaste bakslaget efter upprepade förseningar i NASA:s rymdfärjeprogram . 
Det finns inga planerade uppdrag inför tionde årsdagen av Apollo 11 , och rymdprogrammets framtid är oklar . 
Skylab kommer att störta ner vid en ospecificerad tidpunkt , på en ospecificerad plats . 
NASA beräknar att sannolikheten att en människa träffas av rymdskrot är 1 / 152 . 
Att en stad med minst 100 000 invånare träffas av rymdskrot är en på sju . 
