Jag hade inte kunnat göra detta utan Vox Machina . 
Och inte det som kommer . 
Vad fan hände nyss ? 
Hon tog honom . Raishan tog Thordaks lik . 
Kiki , mår du bra ? 
Såklart jag inte gör . 
Hon gillrade en fälla och vi gick rakt i den . 
Vi visste inte . 
Jag visste . 
Jag har vetat hela tiden , men jag kunde inte övertyga någon . 
Du kan inte beskylla dig själv . 
Det gör jag inte , Vax . 
Varje gång jag tog upp det , varje gång jag höjde rösten , blev jag ifrågasatt , betvivlad , avfärdad . Av min egen grupp . 
Vänta . 
Vad gör du ? 
Jag väntar inte på någons godkännande . 
Jag förlitar mig inte på någon längre . 
- Keyleth , snälla . - Låt bli . Följ inte efter mig . 
Keyleth ! 
Keyleth , hade rätt . 
Vi lurade oss själva . Övertygade varandra att vi kunde lösa allt om vi gjorde det ihop . 
Håller du inte med ? 
Innan Vox Machina var det du och jag . Vi lämnade inget ogjort . 
Du vill ge dig på Ripley . 
Det skulle kännas bra att hämnas mor . 
Det gjorde det inte . För det finns en sak till att ställa till rätta . 
Gruppen då ? 
Det finns ingen grupp längre . 
Om det är det du vill , syster , så stöttar jag dig . 
Vad händer med oss ? 
Fortfarande ingenting ? 
Hans kropp är läkt men han vaknar inte . 
Har du testat att be ? 
Jag vet inte om det hjälper . 
Låt mig prova en sak . 
Scanlan ? 
Hallå , Scanlan ! 
Vakna , ditt lata arsle ! Jag har sprit ! Och nakna kvinnor ! Och nakna kvinnor täckta i sprit ! 
Åh , nej . 
Det fungerar alltid . 
Han kanske inte vill vakna . KAYLIES SÅNG 
Kompis , du kan ha rätt . 
Jag måste hitta Allura . 
Stanna här tills jag kommer tillbaka . 
Okej . 
Förlåt ! Det är Pike , hej . 
Du känner mig . Typ . 
Vilket rum bor Kaylie i ? 
Sex . 
Tack , doktorn . 
Jag är hennes transport . 
Du är helaren . Varför skulle jag kunna göra något ? 
För han bryr sig om dig . På riktigt . 
Jag har inte sett honom känna så för någon annan . 
Jo , sig själv . 
Han har jobbat på en sång . 
Den är till dig . 
Jaså ? 
Varför kom han inte till mig då ? 
Det gjorde han . 
Försökte åtminstone . 
Han riskerade allt för att hitta dig . 
Jag har känt Scanlan länge och vi har varit med om mycket . 
Är ni två , du vet ... 
Nej ! Gud , nej . 
Eller ... Jag menar , okej . 
Jag , du vet ... Vi skulle försöka ... Vi behöver inte prata om det . 
Du får fram något i honom som ingen annan kan och , jag vet inte , du kanske kan få honom att vilja leva . 
Scanlan jävla Shorthalt . 
Så ja , gröna vänner . 
Keyleth . 
Hur ska jag leda asharierna och jag inte kunde få sex personer , sex vänner , att lyssna på mig ? 
Det hör till att göra fel i livet . 
Som mammas trädgård . 
När hon försvann vattnade jag för mycket , för lite ... Allt vissnade . 
Men jag rensade inte bort det . 
Fröna fanns där , precis under ytan , väntade på att komma till liv . 
Fast jag får ingen andra chans . 
Inget spelar någon roll om jag inte hittar Raishan . 
Du vet något . Pappa . Berätta . 
Det finns en gammal ritual . 
Den kan lokalisera någon på stora avstånd . 
Det är precis vad jag behöver . 
Hur använder jag den ? 
Det gör du inte . 
Ritualen är extremt farlig , endast ett fåtal jordashari känner till den . 
De avslöjar den inte utan rådets tillstånd . 
Kalla till ett möte . 
Stilben . Här bor rikets opålitligaste motbjudande människor . 
Är du säker på det här ? 
Men kan inte rensa världen utan att bli smutsig . 
Efter dig , i så fall . 
Korrin , rådet har samlats . 
Vad vill du att vi ska höra ? 
Tack , Uvenda , rådsmedlemmar . Jag ... Det är jag som vill prata med er . 
Jag heter Keyleth , dotter ... Varför är du inte på din aramenté ? 
Jag försäkrar er , vi hade inte kallat er om det inte var brådskande . 
Vid slaget om Emon , stred jag med modiga eldashari som gav sina liv mot Thordak . 
Vi vann . 
Åtminstone tills Raishan förrådde oss . 
Och jag tror ... Jag vet att det är min plikt att stoppa henne . 
Därför ber jag er att anförtro mig jordashariernas lokaliseringsritual . 
Va ? 
Absolut inte . 
Du är inte redo . 
Jag är inte samma tjej som när jag gav mig av . 
Jag har överlevt Feyriket , varit i Avresans helveten . 
Jag har gått igenom eld och blivit ett med den . 
Ni har ingen aning om vad Raishan är kapabel till . 
Ashari har hanterat samma drake förut . 
Våra äldre tillfogade henne en skada som kommer att bli hennes död . 
Vänta . 
Var det vi som gav henne sjukdomen ? Jag visste inte ... Det är mycket som du inte vet , Keyleth . 
Du är inte halvvägs genom dina prövningar . Och nu ber du om vad ? Få hoppa fram i din aramenté och lära dig en farlig rit ? 
Den kan döda dig . 
Jag kan hantera det . 
Kan du ? Det sa din mamma med , och henne har vi inte hört av igen . 
Ashariernas uppgift är att vakta revorna . 
Raishan må beskylla oss för sjukdomen . Du må ha personligt agg mot henne . Men det åsidosätter inte din plikt och det rättfärdigar inte risken . 
Begäran avslås . 
Pappa ? 
Jag är ledsen , Keyleth . 
Jag kan inte lägga mig i beslutet . 
Usla fuskare ! 
Idioter . 
Ni drar till er uppmärksamhet . 
Försvinn ur min åsyn . 
En peppardosa . 
Den här lilla saken . Jag hittade den på Darktowön . 
Du tog fel dörr . 
Jag ville fråga var du fick tag i peppardosan . 
Jag kan svara eller skära halsen av dig . 
Skada inte någon annan som bär mantel . 
Ingen ankarknut i ditt ärr . 
Vi är väl vänner då . 
Vex , lägg av ! 
Syster ! 
Han tänkte döda dig ! 
Nej . Han är med i skrået . 
Ursäkta . Hon är lite ... 
- Hon kan vara lite ... - Oroa dig inte . 
Jag har också en syster . 
Jag älskar henne . 
Ska vi börja om ? 
Du kommer alltid att vara med mig . 
Och en dag är du redo för din egen resa . 
Du måste bara lyssna . 
Ett skepp har tagit sig upp och ner längs Lucidiankusten och levererat dessa vapen . 
Utan flaggor eller symboler . 
Stannar här och fyller på lagret . 
Vet du när skeppet kommer tillbaka ? 
Det kommer bara på natten och meddelar inget i förväg . 
Då får vi sätta oss bekvämt . 
Ni är på egen hand nu . 
Jag beblandar mig inte med de jävlarna . 
Tack , kompis . 
Det finns inga vänner bland tjuvar . 
Kom ihåg , våra skulder betalas med blod . 
Vi ses på andra sidan . 
Må vindarna vaka över er när ni återvänder till era klaner . 
Eldarna släcks och rådet avslutas . 
Inte än . 
Vi är inte klara . 
Ni har inte lyssnat på mig . 
Rådet har bestämt , Keyleth . 
Nej , du gjorde det . 
Inte de . 
Jag har hört att striden inte är värd risken . 
Varnad att vara försiktig . Att vänta ut Raishans sjukdom . Att hålla tyst och fortsätta min aramenté . 
Men det är inte ledarskap , det är feghet . 
Du pratar med en självsäkerhet som du inte har förtjänat . 
Din mor visste om ... Jag är inte min mor . 
Min väg är min egen . 
En riktig ledare är villig att ge upp allt för det hon tror på . 
Det är så jag ska vara när jag sitter i rådet som Stormens röst . 
Ja , ashari har en plikt mot vårt folk . Men vi har även en plikt mot Exandria . 
Vi är faktiskt en del av den här världen , och jag är redo att slåss för den . 
Jag är redo att dö för de jag älskar . 
Du kan neka mig , ledare Uvenda . Men jag lämnar inte arenan om jag inte får samma svar från alla i rådet . 
Eftersom ritualen tillhör mitt folk , måste vår åsikt beaktas . 
Vi är ashari men Keyleth har rätt . 
Vi är även exandrier . 
Det är dags att vi börjar agera som det . 
Pa ' tice , du har ingen koppling till draken . 
Du kan inte utföra ritualen åt henne . 
Därför ska jag lära flickan . 
Instämmer resten av er ? 
Tack för att ni står upp för min dotter . 
Vänta med tacket , Korrin . 
Att få rådets godkännande var lätt jämfört med vad som väntar . 
Många har dött av den här riten . 
När börjar vi ? 
Fortfarande inget . 
Vi borde gå dit och tvinga någon att prata . 
Stubby , jag vet att du vill hitta henne , men vi måste sansa oss . 
Självklart . 
Metodiskt . 
Vad säger du ? 
Jag kollar om jag hör något . 
Du stannar här . 
Toppen . 
Det tar år för jordashari att bemästra sina krafter . 
Att dra energi från marken , bli ett med jorden . 
Men den här platsen , en knutpunkt av korsande mystiska leylinjer , hjälper dig att komma åt samma förmågor . 
Märkliga statyer . 
Ritualen utnyttjar knutpunktens kraft . Men även här är den svår att bemästra . 
Vänta ... Var det här människor ? 
Kom ihåg vad du besitter som ashari . 
Vindens kraft som blåser i ditt hår , stenens kraft under dina fötter . 
Likt leylinjerna , är du en axel som elementen flödar runt . 
Och så snart du har lärt mig , ska jag använda de sakerna . 
Men det kan jag inte . 
För jag har redan förmågan . 
Likt en mäktig alm som gror från ett enda frö , måste du ankra din kraft och låta den växa . 
Ett skepp ! 
Färdigväntat . 
Jag ska inte missa henne . 
Sätt igång ! Ska ske . 
Dålig vana . 
Såna tar död på en . 
Titta vad vi har här . 
Din tur . 
Vi tog en som snokade i hamnen . 
Fan , Vex . 
Knyt an med marken . Stenarna , leran , bristerna . 
Så här ? 
Bra . 
Sjunk in i det nu , men långsamt . 
Om du förlorar kontrollen kan du förlora dig själv . 
Vilken lugnande tanke . 
Jag ... Jag känner något bittert . 
Ja . Fiendeskapets band mellan dig och Raishan . 
Det går genom marken som en sjuk rot . 
Följ det genom jorden . Genom stenen . 
Följ det till henne . 
Ledare ? Det ... Det är för mycket . 
Jag kan inte behålla kontakten . 
Behåll fokuset , Keyleth . 
Nej ! 
Det drar ner mig ! 
Keyleth ? 
Varför klarar jag det inte ? 
Vad fan gör du här ? 
Inget . Jag gick vilse . 
Nu är du upphittad . 
Ledsen , gumman . Lätta ankar . 
Vänta . 
Chefen bad mig att göra det . 
Varför ? Varför bryr hon sig ? 
Vill du fråga henne ? Varsågod . 
Intressant ... Var är din krok , Nikolai ? 
Ja , ja . Jag försökte åtminstone . 
Nej ! Fan ! 
Vad i helvete tänkte du ? 
Du förstörde det nästan ! 
Förlåt . Jag ... Om jag stannar upp ens för ett ögonblick , kommer allt jag känner för Percy tillbaka . 
Som jag sa , jag stöttar dig . Men det fungerar bara om du stöttar mig . 
Jag vet . 
Och det gör jag . 
Hallå ! Inkräktare ! 
Lossa förtöjningen ! 
Sjösätt skeppet ! 
Så gick det med det lugna sättet . 
Vex ! Lite hjälp ! 
Jäklar ! 
Tack , syrran . 
Naturen känner av när något håller dig tillbaka . 
Försök igen . 
Fokusera . 
Knyt an till jorden igen . 
Jag ska inte misslyckas . 
Är det Raishan ? 
Nej . 
Det är något annat . 
Det ser lugnt ut . 
Välkomna ombord . 
Ripley . 
Till er tjänst . 
Fan . 
