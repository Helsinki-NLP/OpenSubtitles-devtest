Pengarna eller livet ! 
Ut ! 
Ut , sa jag ! 
Försiktigt ! Vi vill inte göra damerna upprörda . 
Herregud , nej . 
Vi vill inte skrämma dem - till att berätta var deras smycken ... - Här borta ! Och sånt är gömt . 
Vi vill att de berättar av egen vilja . 
- Definiera vilja , Algernon . - Ursäkta , chefen ? 
Viljans makt att göra saker frivilligt . 
Ni får ursäkta matematikerna . 
Deras huvuden är så fulla av algebra och geometri att de glömmer att uppföra sig . 
Det som händer nu är att Algernon och Chumley går igenom era saker , medan jag underhåller er med min charm - och munterhet . - Chefen , han har en kniv . 
Försök inget med mig , solstråle , för då överlever du inte . 
Okej . 
Händerna . 
Chefen ! 
Vad är det här ? 
Jag tar hand om det . Gå och frikänn dig själv med vördnad . 
Snygga kläder . 
Jag kan se mig själv paradera runt i de stövlarna . 
När du är redo . 
- Du är ... 
- Vad ? 
Inte en man . 
Och ? 
Är det guld ? 
- Är vad guld ? 
- Ringen på ditt finger . 
Åh , ja . 
Jag tror att du kanske måste donera den . 
Jag tror inte att du hörde mig . - Jag sa ... - Jag hörde dig . 
Jag ignorerade dig bara . Ett varningens ord , du vill inte bråka med mig . 
Jag gillar dig . Nej , det gör jag . Du är min typ av kvinna . 
Tyvärr , - måste affärer komma före nöjen . - Okej . 
Gör som du blir tillsagd . 
Kom igen . 
Är ni okej ? 
Hej . 
- Herregud . 
- Vad ? 
Kom igen . Här borta . Sparka den . 
Kom igen . Här . 
Fortsätt . 
Kom igen . 
- Du är okej . - Ta den . 
Förlåt , herrn . 
- Vad är det här ? 
- Grisblåsa . 
Har det hänt nåt här ? 
Thomas Blancheford bråkar . 
Herregud . 
Vem av er är George ? 
Hämta pappa . 
Pappa ! Affären . 
Servera honom , tjejen . 
Du vet var sorbeten bor . 
Hon vill inte ha sorbet . Hon vill ha dig . 
Hon ? 
Hej , pappa . 
Roxy . 
Var är Roxy ? Roxy ! 
- Nell är tillbaka ! 
- Va ? 
Nell ! Din Nell ! Hon är tillbaka . 
Nell är död . 
Jag är änka . 
Kapten Jackson är död . Han dog . 
Han sprängdes itu i slaget vid Blenheim . 
Och du med honom . Det hörde vi . 
Jag undrade varför alla såg så konstigt på mig . 
Saken är den att jag undrar om jag kan bo här i några nätter . 
Jag trodde inte att du ville ha med oss att göra . 
Det var det sista du sa innan du kom in genom dörren med din snofsiga kapten . 
Tja ... Jag har mognat sen dess . Nell ? Nelly ! 
Låt mig se på dig . Se på dig . 
Kalla mig inte Nelly . 
Okej . 
Vad är det här ? 
Pappa betalade inte för en bra . Så vi gjorde den . 
Du retade upp honom när du åkte . 
Får jag dra upp den ? 
Den ger mig kalla kårar . 
Varsågod , Nelly . 
Nell . Förlåt . 
Nu går vi . 
Varför bråkar lord Blancheford ? 
Det är inte lorden . 
- Det är hans son . 
- Thomas . 
- Minns du honom ? 
- Nej . - Han växte upp . 
- Elak och dum . 
Han tycker att det här är kul . 
Varför gör ingen nåt ? 
Vi är hans hyresgäster . 
Eller blir , när nåt händer hans farsa . 
Roxy , alla mina grannar är på krigsstigen . 
Roxanne , bäst att du skyndar dig . 
Kan du säga att min syster är tillbaka från de döda ? 
Det gjorde jag . Hon sa att det inte kan hända . 
- Ohoj , Nelly . 
- Okej . 
- Bäst att jag går . - Ja . 
- Det här är sista varningen . 
- Du måste smöra för pappa . - Det ska jag . 
Det värsta med Thomas är att han är tänd på Roxy . 
- Jaså ? 
- Och han kommer in på värdshuset , full , säger saker , och pappa vågar inte göra nåt . 
Ta hand om min häst , pojk . 
Är du hungrig ? 
" Ja , vi äter hö . " 
Du ska få lite hö . 
Har han slagit dig igen ? 
" Ja , men jag gav igen . Jag kastade av honom , två gånger . " 
Snyggt . 
Herrn . 
God eftermiddag . 
I morse , Thomas , tog min steward emot en delegation från byn med en otrolig historia om att du hade skjutit en mans häst . 
Det var en olycka . 
De sa att du var full , att du red upp och ner för gatan och terroriserade folk . 
Hästen var Nathan Hallidays levebröd . 
Förstår du ingenting om de här människornas liv ? 
Jag är deras rådman . De söker rättvisa från mig . 
En dag , Gud hjälpe dem , kommer de till dig . 
Skrattar du åt mig ? 
Absolut inte . 
Jag drar in din veckopeng . 
- Va ? - Tills den dagen då jag kan lita på att du uppför dig . 
Tvinga mig inte att göra dig arvlös . 
Det är minsann frestande , för din syster skulle vara tusen gånger mer pålitlig . 
Väx upp . 
För Guds skull . För allas skull . 
Håll dig borta från byn tills dess . 
Är det sant att du inte betalade för en riktig gravsten åt mig ? 
Hon kan sova i skjulet med åsnan . 
- Bara en natt . Säg det till henne . 
- En natt ? 
Du krossade mitt hjärta . Du gör det inte två gånger . 
Okej . En natt . 
Okej . 
Du kan bo i huset . 
- Men du jobbar . 
- När gjorde jag inte det ? 
Sätt på dig ordentliga kläder . 
Jag har ingen klänning . 
Titta i skåpet . 
Jag behöll Elizabeths saker . 
Han hade nog köpt en gravsten åt dig . Men jag tror inte att han gillade tanken på dig död . 
Tack . 
Du ser precis ut som din mor . 
Kom hit . 
Ta för er ! Hugg in ! 
Det är inte varje dag en mans dotter kommer tillbaka från de döda ! 
Det är ett mirakel , Sam Trotter ! 
Du , George . 
Hämta Nelly , tjejen . Alla vill ha en glimt . 
Gå nu . 
Hon kommer ner . 
Det ser bra ut . Få se framifrån . 
Du ser så bra ut , Nell . 
- Jaså ? - Ja . Är den bekväm ? 
Nej . Vad handlar det här om ? 
- Saknar du honom ? Kapten Jackson ? - Nell ! 
Pappa vill att du kommer ner nu . 
Alla vill se dig med egna ögon . 
Alla vill höra om kriget . 
Var är ditt svärd ? 
Jag saknar honom lite . 
Förutom ... Jag tror inte att han har lämnat mig , även om han är död . 
Det är som i dag , jag blev rånad av stråtrövare . 
- Nähä ? 
- Och en av dem slog mig . Jo . 
Och det är som ... Jag vet inte , något händer inuti mig . Och ... ni skulle ha sett mig . 
Jag är oåtkomlig . 
Det är han . 
Thomas . 
- Ja ! Buckleigh , din pajas . - Ja . 
Kom hit . 
- Ja . - Ett försprång . 
Kom igen , grabben . 
Firar du något , Trotter ? 
Nej . 
Var är din dotter ? 
- Vilken av dem ? 
- Jag vill träffa henne . 
Jag vill att hon tjänar mig . 
Och Trotter ... Trotter . 
Jag ber dig inte . 
Jag beordrar dig . 
- Jag ska se om jag kan hitta henne . 
- Ja , gör det . 
Vad är det , Halliday ? 
Du ser ut som om din häst har blivit skjuten . 
- Vad är det här ? 
- Det är min äldsta , Nell . 
Hej . Är inte du död ? 
- Var du ute efter nåt ? 
- Jag ville ha den andra . 
Den kommer inte . 
Hon gillar inte dig . 
Hon gillar inte hur du ser på henne eller vad du säger . Och vet du vad ? 
Inte jag heller . 
Jag vill att du går nu . 
Ta dina små idioter med dig . 
Jag ... Tack . 
Hallå där . 
Du kan ha gjort misstaget att anta att jag inte skulle skada en kvinna . 
- Vänta . 
- Men nu vet du bättre . 
- In med dig . 
- Nell . 
Nej ! 
- Nell . - Ta henne ! - Backa ! 
- Slå ner honom . 
- Vart ska du ? - Rör henne inte ! - Nell ? - Du är en stor flicka . 
Sluta ! 
Släpp henne ! 
- Du tvingade mig . - Nell ! 
Du fick mig att göra det här . 
Hon sa att hon var oåtkomlig . 
Nell ! 
Sluta , snälla ! 
- Det räcker ! 
- Sluta . 
Upp med dig , Nell , fort ! Upp med dig ! 
Nell ! 
Spring , Nell ! Spring , fort ! 
- Nell ! 
- Herregud . 
Pappa , säg åt honom ! 
- Herregud . Sluta ! Snälla ! - Låt henne vara ! 
Snälla , sluta ! 
Låt henne vara ! 
Kom igen , Nelly ! 
Kom igen , Nelly . 
- Kom igen , Nell ! - Har du mer ? 
- Ja , Nelly ! - Du då ? 
Ja , Nelly Jackson ! 
- Såg du det ? 
- Vad ? 
Ljuset ? 
Pricken av nåt som svävar ovanför Nells ... Nell ! 
Nelly Jackson ? 
Skrik inte . Du måste titta upp . 
Jag har funderat på det bästa sättet att presentera mig utan att ge dig en chock , Nelly Jackson . 
Det går inte . 
Självklart är det inte nödvändigt att jag presenterar mig . Men i ditt fall , misstänkte jag att det skulle dyka upp förr eller senare . 
Så tre saker . 
Ett , jag är på din sida . Två , den är inte laddad . 
Och tre , den skulle inte ha nån effekt på mig , för jag är icke-kroppslig . 
- Vad menar du med att du är på min sida ? - Se på mig . 
Jag skyddar dig . 
- Varför ? 
- Vem vet ? 
Det här är viktigare . Jag kan bara skydda dig , Nelly Jackson . 
Jag deltar inte i slumpmässiga våldshandlingar . 
- Vad pratar du om ? 
- Som ikväll . 
Va ? 
Han är en översittare . 
Han är en arrogant tölp som gör folk illa . 
- Han startade inget . Det gjorde du . - Han tänkte göra det . 
- Det är inte poängen . - Vänta . 
Menar du att du lät honom slå mig och kunde ha stoppat det ? 
- Jag stoppade det . 
- Inte tidigare ! 
Som när han tryckte ner mitt ansikte i leran . 
Nell , det är jag , George . Är du okej ? 
Vem skickade dig ? 
Var kommer du ifrån ? Se på dig . 
Vad är du klädd som ? 
Nell ? 
Nej , rör dig inte . 
- Okej . - Vänta där . 
Vad heter du ? 
- Har du ett namn ? - Ja . Billy . Billy Blind . 
Vi ses senare . 
Men vänta . 
Tittar du på mig hela tiden ? 
Herregud , tittar du på mig när jag , du vet , - gör det nödvändiga ? - Nell ! 
- Vem pratar du med ? 
- Mig själv . 
- Är du okej ? 
- Ja , jag hörde bara ett ljud , så ... 
Det måste ha varit mössen under golvbrädorna . 
Det var lysande , tidigare . 
Ja , ja . Tack . Ja . - Kan du lära mig hur man ... - Ja . Visst . Kanske . 
Nej . Jag vet inte . 
- God natt . - God natt . God natt . 
Billy ? 
Billy ? 
Billy Blind ! 
Billy ? 
Billy Blind ? 
Poynton . 
Thomas . Kära nån ! Vad gör du här ? 
Jösses . Vilket fult blåmärke . 
Jag åkte hem till dig , men din betjänt sa att du var här . 
- Har du en minut eller två ? 
- Om det är allt . 
Debatten bara fortsatte . Hennes Majestät är så kapabel , till det att hon hör alla sidor . 
Var det hon ? 
Gillar du henne inte ? 
Hur kan jag hjälpa dig ? 
På sistone , har det varit svårt och jag har ingen att prata med , och jag vet att du är upptagen . 
Berätta vad som gör dig upprörd . 
Jag har skulder som min far inte känner till . 
Skulder jag bara kan betala när jag får mitt arv . 
Åtminstone för att han ... dragit in min veckopeng . 
Du sa en gång ... att en man kan sälja sin själ till mörkret . Och i gengäld får han allt han önskar . 
Och att du ... är en person som kan ingripa i sådana frågor . 
Jag vill ha min egendom , Poynton . Jag vill ha allt ... nu . 
Det är ett stort beslut , Thomas . Men om det verkligen är vad du vill , måste du bevisa för mig att du ... har vad som krävs . 
Hur då ? 
Det har inte varit så här städat på åratal . 
Jag kommer aldrig att bli nåt av att bara sitta här . 
Vad hade du tänkt dig ? 
Du gillar det inte . 
Så du tänker ta drottningens shilling ? Hur då ? 
Måste man inte vara soldat ? 
Jag har sett många kvinnor gå med i armén . 
De klär ut sig till män och går ut . Man ser världen , träffar folk och sen ... spränger de dem i luften . 
Skriv den här gången . Så vi vet var du är och att du inte är död . 
Jag kan inte skriva . 
Hitta nån som kan . 
Du kan inte läsa . 
George kan . 
Prästen lärde henne . Hon läser bättre än han . 
Trevligt att träffas , Nelly . Nell . 
Dig med , tjejen . 
Kom , Ashrumbs . 
Hon är åtminstone inte död längre . 
Ja . 
Gå . 
Pappa ? 
Pappa ? 
Jag har skickat skogvaktaren och vaktmästaren till byn med kroppen . 
Jag sa åt dem att säga till hans barn att han blev skjuten under en tjuvjakt . 
Vad höll du på med ? 
Thomas ville skrämmas och lära honom en läxa , vi visste inte ... Vi visste inte att hans hjärta skulle brista . 
Inser du att genom att dölja sanningen gör jag mig själv lika skyldig som du ? 
Jamie , Buckleigh , åk hem . 
Prata aldrig om det här med nån . Då blir du hängd . 
Jag vill aldrig se någon av er igen . 
Ni äcklar mig . 
Förlåt att jag knackar på . Ni känner inte mig , men jag jobbar för lord Blancheford . 
Och ... 
Er far sköts inte vid en tjuvjakt . 
Han blev misshandlad av mäster Thomas och hans vänner . 
De kom hit under natten och tog honom . 
Det gick för långt . Nu försöker de mörklägga det . 
Hur vet du det ? 
Jag hörde skogvaktaren och vaktmästaren prata . 
Lord Blancheford har gett dem pengar för att hålla tyst . 
Jag borde inte berätta det , men jag vet inte . Jag har sett dig i byn ett par gånger ... - Är det din häst ? 
- Åh , nej . 
Jo . Det är en av lord Blanchefords . 
Vad heter du ? 
Rasselas . 
Vart skulle du ta vägen om du tog drottningens shilling ? 
Vems fel är det ? 
Ni vet inte vem jag är . Ni kan inte ... 
- Släpp mig , sa jag ! Släpp ! - Ut ! 
Dumma häxa ! 
Så jag är en kvinna ! Än sen ? 
Jag kan slå ihop era huvuden . 
Förlåt , det var det roligaste jag har sett på hela veckan . 
Jag känner dig . 
Charles Devereux , madam . 
Snobb . Bon viveur . Slöseri med utrymme . 
Men en stor beundrare av skönhet , i vilken form den än väljer att kasta sig upp i . 
Förlåt , jag borde inte ha skrattat . 
Det är så ädelt , att vilja anmäla sig för drottning och fosterland . 
Jag skulle aldrig göra det . Aldrig i livet . 
Jag bryr mig inte om vem som sitter på Spaniens tron . 
Varför skulle jag ? Varför skulle nån av oss ? 
Låt honom hållas , tycker jag . 
Men det är ju trevligt att vara en världsspelare . Kul att fuska lite med grenar . 
Framstegsmarsch , maktbalansen , bla , bla , bla . 
Får jag bjuda på en drink ? 
Du är Isambard Tulley . 
Det hoppas jag verkligen inte . Han har en belöning på 20 pund . 
Ja . 
Amerika , Nell Jackson . 
Den nya världen . 
Det är vad du vill göra . 
Det är du gjord för . Jag känner lukten av det . 
En äventyrlig själ som du , det finns stora förmögenheter att tjäna . 
Herre , ja ! Mahogny , hampa , bomull , tobak . 
Det är vad jag skulle göra om jag var du . Jag kan säga ... Ursäkta , får jag ... ? 
- Pappa är död , Nell . 
- De sa att han sköts under jakten ... - Det är lögn ! 
Mr Rasselas berättade det . 
- Det här är mr Rasselas . 
- Det var Thomas Blancheford . 
- Men hur ? 
- Han kom på natten . Han tog honom . 
Nej , det tillåter jag inte . Han får inte komma undan med det . 
Ta min häst , Nell . Det går fortare . 
Han är ingenting . En nolla . 
Han driver den lokala krogen . 
Jag jagade ut honom ur stan i skydd av mörkret , och sen ... dödade jag honom . 
Utan anledning . 
Bara för att jag kunde . 
Att förgöra en sån man är intressant , Thomas . Men det är knappast något som skapar ett gott rykte . 
Om du vill ha allt nu , om du fortfarande vill det ... Lyssna noga , Thomas . 
- Döda . - Allt du behöver göra är att lyssna . 
Du förstår , Thomas , i det här livet hjälper världen de som hjälper sig själva . Och den här världen behöver män som är kapabla till extraordinära saker . 
Vad står mellan dig och din egendom ? 
Dödade du fel person ? 
Min far . 
Vill du att jag ska döda min egen far ? Nej . Jag vill ingenting . 
Åh , nej . Det är du som vill saker . Och ibland är svaret på ett problem mycket mer prosaiskt och uppenbart än det först verkar . 
Du har rätt . Kulorna gick in efter att han var död . 
Hur vet du det ? 
Jag har lagt om fler sår och lik än du har ätit varma middagar . 
Ingen blodförlust . Hans hjärta hade slutat slå innan de sköt honom . 
Krutet , det gjordes på nära håll . 
Så skjuter man inte tjuvjägare . 
- Vad ska vi göra ? 
- Jag kan inte andas här . 
Jag måste gå . 
Du säger väl inte att jag sa nåt ? 
Tack för att du hjälper oss . 
Det finns ondska i etern , Nelly Jackson . 
- Jag är så ledsen - Det är mitt fel . Om jag inte hade lagt mig i och spöat Thomas . 
Jag måste åka dit - och titta in ... - Gå genom rätta kanaler . 
Va ? Ursäkta , vem är du ? 
Varför är du här ? 
Ni behöver en rådman . 
Lord Blancheford är vår rådman . Han mörklägger det . 
Det blir intressant att höra vad han har att säga . 
- Ge honom ett kryphål . 
- Ett vad ? 
Säg att du misstänker mörkläggning . Men du vet att han aldrig skulle vara inblandad i nåt så tarvligt . 
Se vad som hände när du stormade in . 
- Nej ... 
Om du gör nåt förhastat hjälper jag dig inte . 
Sam Trotters barn är här . De vill träffa dig . 
Jag är ledsen för er far . 
Han var en bra hyresgäst , men han visste vad straffet för ... Min far skulle hellre hugga av sig handen än stjäla från dig . 
- Faktum kvarstår . - Han sköts efter att han var död . 
- Han sköts på nära håll . - Ja , hör på , - du vill inte höra det ... - Din Thomas dödade honom . 
Han och hans dumma vänner och nu försöker du dölja det . 
Inte du . Uppenbarligen . 
Vi vet att du inte skulle blanda dig i något så ... tarvligt . Men någon gjorde det . 
Ni är upprörda , ni låter fantasin skena iväg med er . Men ni uppnår inget genom att hitta på er egen version av händelserna . 
Om jag tvingas hitta en annan rådman , gör jag det . 
Då blir det ditt ord mot mitt . 
Du hördes prata med din skogvaktare . 
Vem hörde det ? 
Du betalade honom och en av dina män för att göra ditt smutsjobb . 
Jag vill erbjuda dig arrendet av Talbot . 
- Va ? - Och i gengäld vill jag inte höra fler vilda anklagelser mot min son . 
Tänk på saken . 
Jag vill inte göra er hemlösa . 
Ingen av er . 
Om vi accepterar det , så accepterar vi lögnen . Att pappa är en tjuvskytt . 
Han skulle inte bry sig om det . 
- Han skulle bry sig om Talbot . 
- De smutskastar honom . 
Talbot är bara en pub . 
Det är vårt hem . 
Det är pappas pub . 
Jag vill inte åka , Nell . 
Okej . 
Verkligen ? 
Vi tar arrendet . 
Armén , då ? 
Det kan vänta tills ni inte behöver mig längre . 
Jag stannar tills dess . 
Halliday ? 
Vad gör du ? 
Jag ska träffa er far , sir . 
Om vad ? 
Arrendet till Talbot . Det kan verka lite förhastat , men om det är ledigt vill jag diskutera villkoren . 
Nej , jag har erbjudit Nell Jackson arrendet . 
Du måste be Halliday att gå . 
- Har hon accepterat det ? 
- Inte än . Jag hoppas att hon gör det när hon är lugnare . För då , Thomas , kanske hon släpper det . 
Jag ska berätta varför . 
De vet . De vet vad som hände . 
Låt dem gå . 
Om det inte har accepterats , låt dem gå . Det är bättre så här . 
Halliday är pålitlig . Han vet vad han gör . 
Sen när är du intresserad av att främja en god mans sak ? 
Jag har varit ovärdig dig . 
Jag har förödmjukat dig och låtit mig påverkas av fel människor . 
Och jag är ledsen . 
Jag vill lägga det bakom mig ... Så det räcker inte att göra dem föräldralösa . Ska du göra dem hemlösa också ? 
Säg inte så . 
Ur syn , ur sinn . 
Det är frestande . 
De är unga och starka . 
De hittar andra vägar att följa . 
- Vad är det ? - Jag företräder lord Blancheford . Här är er uppsägning . 
Vad pratar du om ? Han erbjöd mig arrendet i går . 
Ni har till kl. 12 på er att packa . 
- 12 ? - Är du dum ? 
- Han erbjöd mig arrendet ! 
- Allt som är kvar sen - rensar jag ut åt er . - Jaså ? 
Jag skulle börja packa . 
- Vad ska vi göra ? 
- Jag vet vad jag ska göra . 
Vad ? 
- Ur vägen ! Var är han ? - Du kan inte gå in , kom tillbaka ! 
Jag vill prata med dig . 
Jag kunde inte stoppa henne . 
Ingen fara , mrs Belgrave . 
Jag har inte hört av dig . 
- Jag antog att du inte ville ha arrendet . 
- Lögnare . 
Du kommer undan med allt , eller hur ? 
Till och med mord . 
Din far åkte fast för tjuvjakt . 
Sluta säga så . Vi vet alla att det inte är sant . 
Du kommer troligen undan med det . Mörda min far och märka honom som en brottsling . Den ärligaste mannen någonsin , bara för att dölja vad tölpen gjort . 
Jag vet att du kommer undan med det , såna som ni gör alltid det . Men du förstår väl om jag är lite upprörd ? 
Vad kan jag göra för att övertala dig att lägga ner den där ? 
Okej . 
Jag ger dig arrendet . Jag ger dig vad som helst , tio pund , 20 . 
Du kan inte lita på henne . 
Skulle hon går härifrån utan att berätta att du mutat henne ? 
Skulle jag ta emot pengar för att hålla tyst om att den här värdelösa bandhögen dödade min far ? 
- Jag tror inte det . 
- Din idiot . 
Jag var en idiot som försökte skydda dig . 
- Du ska ställas inför rätta . - Nej . Va ? Nej ! 
Jag tänker inte dras ner och förödmjukas av dig längre . 
Du ska ta konsekvenserna av det du har gjort . Nej ! 
Den var inte laddad . 
Den här är det . 
Kom igen då . 
Gör ett försök . 
Se vad det gör för nytta . 
Nej . 
Din djävul . Din fasa . 
Din fördömda präst från helvetet . 
Hon dödade honom ! 
Hon sköt honom ! 
Hon mördade min far ! Mord ! 
- Mord ! - Lögnare ! 
Du är en lögnare . 
Det var du som kom hit beväpnad och hotfull . Nu har du en tom pistol i fickan . 
Ur vägen . 
Du hängs för det här . 
Det tänker jag inte göra . 
Hon såg vad som hände . Du såg vad som hände , Sofia . 
Du såg vad som hände . 
- Du berättar sanningen . 
- Hon mördade lord Blancheford ! 
Nej , det gjorde jag inte ! 
Det var han . 
Nej , det var han . Det var han . Han dödade sin egen far ! 
Rasselas , jag gjorde det inte . Tror du mig ? 
Tror du mig ? 
- Du tror mig , kom igen . 
- Gör nåt . 
Vad händer ? 
Stoppa henne . 
Släpp mig . 
Snälla . 
Efter henne ! 
Hon säger att hon inte gjorde det . 
Vem gjorde det ? 
Sofia ? 
Det var hon . 
Jag tror dig inte . 
Vad gör du ? 
Rasselas ! 
Ta en av hästarna och hämta en rådman ! 
Fort ! 
George , Roxy , kom ut hit nu ! 
- Roxy ! 
- George , Roxy ! Kom ut hit nu , vi ska åka ! 
- Vad händer ? 
- Kom igen . 
- Vi behöver våra saker . - Glöm dem . Nu , sa jag ! 
Kom igen , fort . 
- Skynda på ! Rasselas , nu ! - Roxy , kom igen . Upp med dig . Kom igen , Roxy . 
