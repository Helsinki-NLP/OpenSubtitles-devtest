Ray , Ray ? Hur är det ? Hallå ? - Jag är hans fru . 
- Ring efter ambulans , nån ! Har ni ringt ambulans ? 
- Ojämn puls . - Intravenöst i höger arm . 
Okej . Se till att hans syrenivå är åtta liter . 
Han behöver EKG , full blodstatus och transfusionsstatus . 
Han har hjärtflimmer , kolla pulsen . 
Ingen puls . 
- Hej , raring . 
- Jag är hemma med barnen . Hur mår han ? 
Han opereras nu . - Då Raymond Horgan ... - Okej . - Jag håller dig underrättad . - Okej . - Jag älskar dig . - Hej då . ... efter att ha drabbats av en hjärtinfarkt . - Absolut en oväntad händelseutveckling . - Jösses . Vi vet inte om rättegången kommer att fortsätta just nu . 
Rae , finns det nåt prejudikat för att sånt här händer ? En svaranden som hoppar in och räddar sin advokats liv ? 
Det brukar faktiskt vara tvärtom . Men som svar på frågan finns ingen regel . Det är upp till domaren . 
Och med tanke på domaren här , vet man aldrig . 
Om rättegången ogiltigförklaras , börjar man om från noll ? Det verkar så . 
Det här är åt helvete . 
Vill du ha nåt att dricka ? Lite vatten eller nånting ? 
Ja . - Ja , tack . - Ja ? 
Lorraine , jag vill bara beklaga . Och om jag kan hjälpa ... Det låter väl ihåligt , men om jag kan göra nåt ... 
- Tack . - Okej . - Okej . - Tack . 
- Mrs Horgan ? - Ja ? - Mrs Horgan ? 
- Ja . Han kommer att klara sig . Och kanske må ännu bättre . 
- Säkert ? - Det var ingen hjärtinfarkt . - Det var bradykardi . - Åh ... Ett elektriskt problem som saktade ner hans hjärtrytm till nära noll . Vi satte in en pacemaker . Ingen neurologisk skada . 
- Han går härifrån piggare . - Tack , doktorn . 
Så han blir bra ? 
- Han kommer att bli bra . - Ja . Bättre . Han är i uppvakningen nu . 
Om några timmar är han på salen , och då kan du träffa honom . Åh , herregud . 
- Tack . - Ingen orsak . Ja ? 
Vi har ett problem . 
Ja , vi har ett problem . 
Juryn såg just Rusty uppträda osjälviskt och ... Vi måste få rättegången ogiltigförklarad . - Va ? - Ja . - Vi ... - Vi vinner ju . 
- Jag undrar det . 
- Ogiltigförklarad rättegång , han går fri . - Nej . Det vet vi inte . 
- Jo , det gör vi . Kom igen . Andra gången lär han veta vår plan . Tänk efter lite . För att vara en lögnaktig psykopat - är han rätt charmig , visst ? - Det är ... Och han räddade nyss ett människoliv inför juryn . Det kan också hävdas att juryn såg honom agera impulsivt , på samma sätt som han gick överstyr . Men man måste lita på juryn . 
De är bättre utrustade att visualisera händelserna den kvällen än nån av oss två . 
Frågan är vad som händer nu . 
Man kan inte fortsätta utan huvudadvokat så långt in i en mordrättegång . 
De kanske pausar allting ? 
Jag tror inte att det funkar så . 
Av allt juridikexperterna säger , så ... Så , vad tänker vi ? 
Tänker vi ? 
Mr Delay Guardia , du är väldigt förtegen av dig . 
Jag sitter och väger principerna om rättegångsekonomi mot dito om rättvisa . Som rättens ombud inser vi att vi har en plikt att tillse att rättegångar är fria från fördomar och partiskhet . Vad i helvete pratar du om ? Det var länge sen vi läste juridik . 
- Vad pratar du om ? - Jag menar att vi anser att rättegången bör ogiltigförklaras . 
- Det hade räckt att säga det . - Vi säger nej . 
Vill ni fortsätta ? 
Jag är beredd att ta över . 
- Genast ? 
- Ska du ta över ? 
Imorgon . Jag behöver en dag . 
Mr Delay Guardia ? 
Förlåt . Jadå . Åklagarsidan är redo att fortsätta . 
Jag vill företräda mig själv . 
Ursäkta ? 
Jag vill ta över som förstaadvokat . Jag är redan inne i fallet och har mer erfarenhet än ms Winslow . - Man kan inte vara vittne ... - Hon kan biträda mig . ... och advokat i samma rättegång . Jag kommer inte att vittna . Det slår jag fast . Du kommer att vittna och vara tidernas slugaste vittne , för du kan lägga fram din sak för juryn och påverka dem ... 
- Min advokat är sjuk . - ... men slippa korsförhör . Jag ska inte vittna till min egen fördel . Jag påminner domaren om att detta är min rätt . 
Då får jag i min tur påminna dig , mr Sabich . Vid minsta antydan att ge din version av kvällen låter jag åklagarsidan sätta dig i vittnesbåset , där du kommer att bli korsförhörd fullt ut . 
Och om du skjuter dig i foten , kan du inte överklaga grundat på sjätte tillägget att ha en inkompetent advokat . 
Tänker du företräda dig själv ? 
Så länge han inte vittnar finns det inget som hindrar . 
Jag förstår , fru ordförande . 
Dålig idé . Men du får skylla dig själv . 
Jag ska instruera juryn , och vi fortsätter imorgon kl 10 : 00 . 
Du har tid att ändra dig . 
Hur är det möjligt ? Ni lovade att skydda honom . 
- Vi ska göra vårt bästa . - Ert bästa ? Ni ska göra ert bästa ? 
Har ingen omsorg om min son ? 
Han ska nu korsförhöras av mannen som mördade hans mor . 
- Han har rätt att representera ... 
- Han är en mördare ! 
Det här är ett fall med många vändningar , men detta är ändå en sensation . 
Eleanor , detta med att Rusty Sabich företräder sig själv , - vad tänker du ? - Mamma , det här är galet . 
Underskatta inte din pappa , vännen . - Inte som jurist . 
- Mamma , kom igen . Det är fan sjukt . 
Sluta ! Sluta . 
Okej , vi ses där inne . 
Ursäkta att jag är sen , fru ordförande . 
Mr Sabich . 
Hej , Michael . Låt mig först framföra mitt djupa deltagande . Jag kan inte föreställa mig smärtan att mista sin mor . 
Du dödade min mor . 
Brukade du åka ofta till din mors hus och bara titta ? 
För att se hennes liv . Att se det liv hon inte ville att du skulle vara en del av . Ja . Sa hon nånsin varför hon inte ville att du skulle vara det ? 
Nej . Berättade din far nånsin varför hon inte ville det ? 
Det måste ha gjort dig ganska arg . 
Kan man uttrycka det så ? 
Inte nog för att döda . Försiktigt . 
- Raymond . 
- Jag bara tittar på . 
Det var intressant , Michael , för de sista veckorna av hennes liv hade du flera sms-växlingar med din mor . 
Skrev du till henne : " Det vore enklare om du var död " ? Sms:ade du det ? 
Hon sårade inte bara mig . Hon sårade min far . " Jag är jävligt arg på dig . Du har förstört mitt liv . " 
Sms:ade du det ? 
Du ville att hon skulle dö . 
Nej , jag sa att det vore enklare . 
Folk går vidare efter dödsfall . Skilsmässa är svårare . Det var det jag menade . 
Okej . Det räcker så . 
Bra . Du filmade mig när jag gick in i din mors hus kvällen hon dog , och du vittnade om att du sett mig gå in där förut . Så du visste att din mor och jag hade en affär . 
Ja . Att hon inte vill ha dig i sitt liv men hade känslor för mig , fick det dig inte att hata mig ? 
Jag hatar dig för att du dödade henne . 
Varsamt , Rusty . 
Efter att du filmat mig , vad gjorde du ? 
Jag stack . Efter att ha sett mig gå in , hur snart gick du därifrån ? 
- Nästan direkt . 
- Vart tog du vägen ? Jag åkte hem . 
Vem var hemma ? Min far . 
Bara ni två ? 
Ja . Nån mer ? 
Nej , bara vi . 
Så ingen kan ge dig alibi utom han . Och bara du kan ge honom alibi . 
- Protest . 
- Avslås . 
Sa du till din far att du sett din mors älskare gå in i hennes hus ? 
Svara på frågan , Michael . 
Jag minns inte om jag sa nåt alls . 
Så är det möjligt ... Är det möjligt att du sa till din far att du såg din mors älskare gå in i hennes hus kvällen hon mördades ? 
Jag minns inte att jag sa nåt alls . 
Ett antal dokument i din dator konfiskerades av polisen . De visade att du hade stort intresse för din mors tidigare fall . 
Du gick ut på sajter om sanna brott och sökte efter information som inte fanns i gängse massmedia , även om Bunny Davis . - Protest . 
- Bifalles . Ställ frågor , advokaten . Han måste passa sig . 
- Dödade du din mor ? - Protest ! Eller din far ? Dödade han din mor ? - Oj . - Säg att du har fog för de frågorna . 
Jag har varken grund för att anklaga vittnet eller hans far . Hur skulle jag kunna det ? Efter en kort och slarvig utredning utförd av polisen , avfördes de från utredningen av åklagaren ... 
- Han går för ... - Domare ! 
Jag frågar , dödade du din mor ? Din sjuka fan ! 
Pappa ! 
- Det räcker ! - Mr Caldwell , kliv tillbaka . 
Vad fan håller ni på med ? 
- Backa . - Kliv tillbaka , mr Caldwell . 
Ni skulle ta hand om honom . 
Mr Sabich , var du rädd när Dalton Caldwell attackerade dig ? 
Raymond hade ett uttryck för när ett fall gick fel , att det var åt skogen , åt helvete , eller åt helvete med besked . 
Det här är nog åt helvete med besked . 
Han framstod desperat . Han anklagar alla utom sig själv . Okej . Okej . Lugn . 
Så han klarlade att nån var där , som bar på hat mot Carolyn Polhemus och som kan ha känt till detaljer om Bunny Davis fall . 
De pekade på Liam Reynolds , och sen pappan som framstod som helt jävla galen . 
Så vi ... Rigo . - Vi kallar Rigo . - Rigo ? - Nej , Rigo är helt på Dustys sida . - Ja . Liksom Eugenia . Ställ rätt frågor . 
- Rigo avskyr mig . - Men inte mig . 
Jag ställer frågorna . - Nej . - Jo . - Jo . - Nej . Jag ska tala om varför . För om vi inte gör det , går vårt fall åt helvete med besked , bortom rimligt tvivel . 
- Vad kommer Rigo att säga ? 
- Jag vet inte . 
Lägg av . Skitsnack . Ni två är vänner . - Säg bara vad hon ... - Nej , ni två är vänner . 
Vad ska hon vittna om ? 
Troligen om det jag såg , Rusty , och det jag ser just nu . 
Vad menar du ? Att du gick helt överstyr , som du gör här och nu . 
Va ... Du vet att jag inte ville vittna , visst ? 
Jag vet att du vet det . 
Har jag fattat helt fel ? 
- Har jag fattat ... - Vad ... Carolyn var en drog . Du var en missbrukare . Missbruk förstör liv . 
Herregud . Det var en sak att förstöra dig , men du tänkte inte låta henne förstöra din familj . 
Herregud . ... att hon tänkte behålla barnet , eller hur ? 
Sa hon den kvällen att hon tänkte behålla barnet ? 
Hon tänkte behålla barnet . - Ditt barn . - Ut ur bilen . 
Ut ur bilen . 
Liam Reynolds var inte inblandad i mordet på Carolyn , men ändå åkte ni två till fängelset för att träffa honom . - Stämmer det ? 
Varför ? 
Vi låter Rusty ge svaret . 
Även om du lät döda Carolyn , kan det bli till din fördel . 
Du måste ha en medbrottsling , alltså hade du nåt att köpslå med . Okej , tänk dig , du avtjänar nu livstid för mordet på Bunny Davis . Men genom att visa oss på Carolyn kan du möjligen bli frigiven . Även om du var inblandad i mordet . 
Nu snackar vi verkligen perverst . 
Bara så att jag förstår , om jag erkänner nåt i en ... - Med medbrottsling . - ... åklagares mord , - kan jag bli frigiven ? - Ja . 
Säkert är att du för närvarande avtjänar livstid utan chans till villkorligt . Jag erbjuder dig en chans att ändra på det . 
Det här är härligt . Nej ! För i jösse namn . 
Jag ... Jag hade ingen jävla aning . 
Du är desperat . 
Förkortat straff i utbyte mot erkännande i mordet på Carolyn Polhemus . 
Jag var inte där . Jag visste inte att han skulle göra så . 
Tog du avstånd från mutförsöket ? Protest ! 
- Bifalles . - Förlåt . Tog du avstånd från denna metod ? 
Ja . När han berättade , sa jag att han hade gått över gränsen . 
Svarade han ? 
Ja , han sa nåt i stil med ... Det gäller mitt liv . Jag gör vadhelst jag måste . 
Vilken hjälte . När du först gavs fallet av svaranden , fick du några särskilda instruktioner angående bevismaterial ? 
Allt bevismaterial , även rättstekniskt , skulle överlämnas enbart till honom . 
Fick du några särskilda instruktioner om vem bevismaterialet , även rättstekniskt , särskilt skulle undanhållas från ? 
Mr Molto och dig . 
Vilken besvikelse . 
Ert vittne . 
Då var det dags . 
Jag försökte desperat bevisa min oskuld , hela tiden , mot anklagelser mot mig som jag ansåg felaktiga . Kan man uttrycka det så ? Okej . Och jag vidhöll hela tiden min oskuld i mordet av Carolyn Polhemus . 
- Eller hur ? 
Enligt din erfarenhet , kriminalinspektör , är det ovanligt att en åklagare ber dig hålla information er emellan ? 
Det är inte ovanligt , nej . 
Och du vet att jag bad dig hålla bevismaterialet mellan oss just därför att jag inte litade på att mr Molto och mr Della Guardia skulle driva en opartisk utredning . Är det en rättvis beskrivning ? 
Tack . 
Hur mår du ? 
Tja , du vet , de ... De kallade två vittnen för att fastställa min ... Jag var lite för ivrig i att bedyra min oskuld . 
Strunt samma . Läget är ändå bra . Vi klarar oss . Har du börjat ta de här igen ? 
Jag behöver fokusera . 
Hur ska jag klara det ? 
Du borde ha talat om det för mig , Rusty . 
- Jättebra . Ja . - Ja . Tack . 
Alla reser sig . 
Rättegången fortsätter . Domare Lyttle leder förhandlingarna . Varsågoda och sitt . 
Jaha , mr Molto . Har åklagarsidan nåt mer ? 
Ja , fru ordförande . 
Åklagarsidan kallar Rusty Sabich . 
Vad fan var det där ? 
Eftersom mr Sabich insisterade på att vittna genom inspektör Rodriguez är det inte mer än rätt att vi får korsförhöra . 
Jag hörde ingen protest . 
Jag såg inget behov , eftersom rätten gjorde det klart att om svaranden antyder en egen version ... Jag vittnade inte . Jag korsförhörde ert vittne . 
Men du bröt mot direktiven . Du vidhöll din oskuld . 
Du kallade vittnet och kriminalinspektören för att påvisa min skuld och ohederlighet . Mina frågor visade min ärlighet och oskuld , helt enligt riktlinjerna . 
Du gav din version . 
Jag varnade dig för att ens introducera ett uns av nåt utanför bevismaterialet ... Och det gjorde du . 
Okej , du har två alternativ . 
Ogiltigförklarad rättegång ? Det får du . Helt enligt reglerna . 
Jag tvingar dig inte att fortsätta . Men om du fortsätter måste du vittna . 
Du öppnade dörren för det här . 
Ta ogiltigförklarad rättegång . 
Jag ska vittna . 
- De ville ha ogiltigförklarad rättegång . - Vad fan ? - Nej . - De höll på att förlora . - Därför kallade de mig ? - Kanske det . Eller så ville de få dig i vittnesbåset där du är ett enkelt mål . 
Okej , sätt mig i vittnesbåset . Okej . Låt Moltos narcissism - bli tydlig för alla . - Varför ? Och din , då ? Vad menar du med det ? 
Gjorde du det med flit ? 
Vadå ? 
- Tror ... - Du introducerade vittnesmål . - Var det medvetet ? - Nej ... Varför skulle jag göra det ? 
För du är Rusty Sabich , och du kan göra vad du vill . 
Mya , kanske , bara kanske gjorde jag det för att jag kan min sak . 
Det tror jag inte . 
Jag hoppar av . 
Rusty Sabich väntas vittna till sitt eget försvar , så han är inte bara svaranden utan sin egen försvarsadvokat . Och han ska även vittna . Va ? 
Han kommer inte att ha ett biträde , vilket betyder att han kommer att köra solo . 
Mycket vilar på hans axlar i den här rättegången . Sabich verkar ha målat in sig i ett hörn . Jag vet inte om nåt annat än ett under ... Herregud , Rusty . ... kan rädda honom ur knipan . 
Piller . Vad för piller ? 
- Han tar Ritalin . 
- Skojar du ? Jag hörde mamma i telefon med sin terapeut . Han brukar visst ta det inför stora rättegångar . 
För att fokusera bättre . Ja . 
Så han tar det innan han vittnar imorgon ? 
Ja , jävligt dumt . 
Är det möjligt att få lite sånt där Rusty Sabich-älvstoft ? 
Jag vet inte om det är nåt jag kan ge dig . 
Säg att du inte har sovit här i natt . 
Nej , jag kom tidigt . 
Okej . Är du redo ? 
Ja , jag är redo . 
Bra . En stor dag . 
Jag tänkte på juristlinjen och hur hårt vi pluggade . 
Ja , ge mig en dag bara , Nico , då jag kan säga att det var värt allt . 
Idag är den dagen , Tommy . 
Det är typ Crime Junkie 101 . Man vittnar inte till sitt eget försvar . 
Men han gjorde ju det . Åklagarsidan kallade honom ... Hur företräder man sig själv utan att verka schizofren ? 
Nåt som kan skapa tvivel hos juryn . 
Hej , Mya . 
Lycka till idag . Jag vill bara säga att nyckeln är att inte låta honom få dig ur balans , vilket är hans avsikt . 
Att provocera dig . Nappa inte på betet . 
Tack , Mya . 
Får jag ge mer allmänna råd ? 
Får jag be om ursäkt först ? 
Ursäkten godtas . 
Du kanske har rätt . 
Jag har jämt rätt . 
Låt honom inte göra dig till en skitstövel . 
Det är inte bra om juryn uppfattar dig så . 
Gör inga medgivanden . 
- Jag kommer att vara där . 
- Nån kom . - Jag måste lägga på . - Okej . 
- Vad gör du här ? 
- Jag är utskriven . 
Du behöver mig . 
Är det verkligen bra för dig att vara i rättssalen ? 
Jadå . Jag är okej , säger läkarna . Och du ? 
Svär du att säga sanningen , hela sanningen och inget annat än sanningen ? - Ja . 
- Varsågod och sitt . 
Mr Sabich du sa att du vidhöll din oskuld hela tiden inför inspektör Rodriguez . 
- Det stämmer . 
- Talade du sanning ? 
Ja . Var du helt sanningsenlig mot henne ? 
Jag avslöjade inte min relation med offret . 
Avslöjade du för henne att du var i offrets hus kvällen för mordet ? 
- Så småningom . - Så småningom ? 
Så när du först tilldelade inspektör Rodriguez fallet i din egenskap av vice chefsåklagare , berättade du att du var på platsen kvällen för mordet ? 
Nej . Berättade du för nån med koppling till fallet ? 
Jag dödade henne inte . 
Är de första 48 timmarna viktigast i varje polisutredning ? 
Och hade det varit till hjälp för polisen och utredarteamet att få veta att du var på platsen ? 
Din poäng är gjord . 
Jag avslöjade inte min närvaro . 
- Var du förälskad i henne ? - Jag blev det . 
Kan man säga att du var fixerad vid henne ? 
Jag var förälskad i henne . Var gränsen går för fixering ... Att skicka 30 sms eller mejl på eller nära dagen för mordet . - Är det fixering ? - Jag var förälskad . 
Kvällen för hennes död , åkte du dit i hoppet att hon skulle ta dig tillbaka ? 
Det stämmer . 
Skickade du följande sms timmarna före hennes död ? 
" Det här är fel . Du kan inte göra så . 
Du får inte behandla mig så här . Svara när jag ringer , för fan . " 
- Skickade du dessa ? - Ja . Och det här ? " Jag vill vara med dig resten av livet . " 
Skrev du detta till Carolyn ? Att du ville vara med henne resten av livet ? 
Jag var kär i henne . 
- Var du arg på henne ? 
- Jag var frustrerad . 
Frustrerad , som i detta sms ? 
" Svara när jag ringer , för fan . Vem fan tror du att du är som behandlar mig så ? " 
Är det frustration , eller kan man kalla det ilska ? 
Jag skulle kalla det passion . 
Passion kan förblinda en . Jag tappade verkligen bort det som är viktigast i mitt liv . Min fru och mina barn . 
Passion är en farlig drog . Du är inte heller immun mot den , Tommy . 
Du är så uppfylld av att få mig fälld att du inte inser faktum att du saknar verkliga bevis . 
Ja , jag var förälskad i henne . Ja , jag avslöjade inte min närvaro , men jag dödade henne inte . 
- Slog du henne med en eldgaffel ? - Jag slog henne aldrig . 
Jag är ingen våldsam person . 
Mr Ratzer , kan du resa dig ? 
Har du mött den personen förut ? 
Det finns en förklaring . 
Här är bilder tagna från ert grannhus . 
Det är ni två , eller hur ? 
Fångar det situationen på ett korrekt sätt ? 
Ordförande , en orättvis överraskning . 
Som genmäle . Vittnet sa nyss att han inte är våldsam av sig . 
Fortsätt . 
Han kom hem till mig oinbjuden . 
Han gjorde intrång och skrämde mig . 
Så du klådde upp honom ? 
Jag är skyldig till att ha handlat i desperation . 
Det fick mig att dölja min relation med Carolyn Polhemus . Det fick mig att ivrigt försöka få ett erkännande från Reynolds angående mordet , och reagera våldsamt mot Brian Ratzer . Förresten kom han till mitt hus och bultade våldsamt på dörren när min dotter öppnade . 
Är jag lättretlig ? Ja , det är jag . 
En person jag älskade mördades brutalt . Jag är anklagad för det brottet . 
Såna omständigheter kan locka fram många saker hos en person , bland annat desperation . Svaghet , känslomässig instabilitet . Jag ber om ursäkt för allt det . 
Jag är skyldig till allt detta . Men jag är inte skyldig till mordet på Carolyn Polhemus . 
Jag tog inte hennes liv . 
Jaha . Och dr Kumagai ? 
Har du nånsin tagit strypgrepp på vår rättsläkare ? 
- Ska jag upprepa frågan ? 
- Nej , jag hörde . Jag fick veta att han hade dolt bevis i ett annat fall . Eller åtminstone underlåtit att ge mig tillgång till det . Stämningen blev upprörd mellan oss och ... Beklagligt nog blev jag våldsam . 
Beklagligt nog tog du stryptag . Nej , det gjorde jag inte . När känslorna kokade - och du grep hans strupe ... - Hans rockslag . Okej , när känslorna kokade och du grep hans rockslag , beslöt du att göra det eller förlorade du kontrollen ? 
Jag vet inte vad frågan var . 
Beslöt du att göra det eller förlorade du kontrollen ? 
Eller mr Ratzer , när du slog honom upprepade gånger som vi såg . Beslöt du det eller förlorade du kontrollen ? 
Han vägrade gå därifrån . 
Vad skulle du göra ? 
Så du förlorade kontrollen . 
Du , se på mig . Se på mig . 
Det där var utomordentligt . 
Det här är rena tortyren . 
Rena tortyren . 
Jag ljuger för min familj hela dagarna . 
När jag är med dem vill jag bara vara med dig . 
Resten av livet , va ? 
Jag minns inte att jag skrev det . Bara nåt man säger ? 
Vad händer nu , om jag vågar fråga ? 
