- MoviesMod.lol Statistik visar att OS-medaljörer följer tre regler inför tävlingar . 
Var utsövd ... Var förberedd ... Och undvik alla distraktioner . 
Här har de utbildats , Nobelpristagare och statsöverhuvuden , författare och vetenskapsmän . 
Och jag kan bli en av dem . 
Där inne väntar min framtid . 
Jag har väntat i åratal . 
Nu är det dags . 
- Hejsan . - Hej . 
- Hej . - Hejsan . 
- Och det här är ... - Jude . 
Ruby . 
- Hej . - Lin , hej . 
Maxton Hall THE WORLD BETWEEN US 
EFTER ROMANEN " SAVE ME " AV MONA KASTEN 
- Hoppas jag inte gör nåt fel . - Inte då . Professorn tar in dig vad du än gör . 
Hade inte din mamma honom som lärare ? 
Lite får vi nog anstränga oss . 
Ja , det får vi nog . Upp med hakan ! 
Alistair ! Vänta ! 
Redo ? 
Självklart . 
Vi behöver bara gå in och få besked att vi har kommit in . 
Ni som inte känner mig , jag heter Jude och går andra året på St Hildas , och jag ska hjälpa er med ansökningen . 
I den första intervjun vill lärarna testa ert kritiska tänkande och om ni kan diskutera ett ämne . 
I den andra , vill de se hur ni arbetar under press . 
Den tredje och sista intervjun handlar om er själva . 
Passar ni in på Oxford ? 
Den är viktigast . 
Första omgången börjar om 45 minuter . Ni hinner gå igenom era anteckningar , kanske äta nåt . 
Ni har kommit så här långt . Oxford vill ha er . 
Försök att inte förstöra för er själva . 
Jag ropar upp er . 
Ruby Bell . St Hildas . 
Lycka till . 
Var inte nervös . Du fixar det . 
Var du nervös ? 
Ja , tio gånger värre än du . 
Men jag kom in . 
Vi ses senare . 
Tack . 
Vi är glada att ni tackade ja till vår inbjudan . 
Tack , så roligt att höra . 
Underbart . Då börjar vi . 
För några år sen publicerade New York Times en debattartikel som hävdade att den brittiska monarkin var en slösaktig anakronism . 
Kan vårt dubbla system med monarki och parlamentarisk demokrati fortleva , eller bör vi bli republik ? 
Frågan kan diskuteras på två sätt . 
Å ena sidan kan man hävda att monarkin ger stabilitet , åtminstone symboliskt . 
Å andra sidan , de enorma kostnader som denna symbol för med sig kan ifrågasättas . Med tanke på alla länder som blomstrar med andra styrelseformer . 
Bra . Fortsätt . 
Marknaden bygger på spekulation , eftersom framtiden tyvärr inte är särskilt förutsägbar . 
Men vinst skapas i nuet , vilket en framgångsrik affärsmodell drar nytta av . 
Tack , mr Beaufort . 
Äpplet faller inte långt från trädet . 
Er far var etta i sin avgångsklass på Balliol . 
Han var ljusår före alla andra med sina kunskaper och sin ambition . 
- Hur gick det ? 
- Du först . 
Bra , tror jag . 
Det var riktigt roligt . 
Jag citerade Platon ... 
De stirrade åtminstone inte på dig . 
Min lärare hade sammanväxta ögonbryn och såg ut som en arg mr Bean . 
Jag tittade på dem hela tiden . 
- Det såg han . - Nej . Hallå . 
Hur var det ? Okej ? 
- Bra . - Ja . 
Ni kan behöva koppla av ikväll . 
I kväll kl. 20.00 ? Oxford-stil ? 
Ja ! 
Här har vi den världsberömda Turf Tavern . 
En pub som har besökts av Liz , Oscar och så Järnladyn själv när hon gick här . 
Där finns det plats . Kom . 
Vem har vi här ? 
Det verkar vara nåt . 
Där är de . 
En specialitet . Ett måste för alla Oxford-besökare . 
Cross Keys . 
Så ser jag också ut när jag dricker vatten . 
Smaka på den här . 18-årig whisky . 
Vad är det för fel ? 
Och bartendrarna måste skriva under ett sekretessavtal för att jobba här . 
Seriöst ? 
Den minen gjorde jag också först . Men senare sprang jag halvnaken över campus och citerade poesi . 
Jag skippar gärna det . 
Då får det vänta tills du är student här . Skål . 
Herregud ! 
Väldigt starkt . 
Jag ska ta lite luft . Min väska ? 
- Aj ! - Du är för uppenbar . 
Ska du säga ? 
Är allt okej ? 
Är frågan retorisk ? 
Är du nervös för intervjuerna ? 
De spelar ingen roll . Jag kan ändå inte börja på Oxford . 
Varför inte ? 
Du har ju varit bäst i klassen två gånger . 
- Om du ... - Jag har gått två månader över tiden . 
Det vore vanvett att behålla det . 
Men jag älskar honom verkligen . 
Och bebisen också . 
Jävla hormoner . 
Det finns studieprogram för mammor . 
Jag såg det när jag letade stipendier . 
Jacinda Ardern fick barn när hon var premiärminister . 
Vi känner inte varann men jag ser ju dig . 
Hur du har kämpat på under ... 
Om nån kan klara det , så är det du . 
Jag fattar varför han inte kan glömma dig . 
Du får allt att verka möjligt . 
Oavsett hur hemskt allt är . 
Vad menar du ? 
Vet du inte hur ledsen han är ? 
Han gjorde ju slut . 
Ibland visar man sin kärlek genom att släppa den . 
OS-poäng efter en dag i Oxford : 
Sömn : noll . Distraktion : tio . 
Bra jobbat , Ruby Bell . 
Du imponerade på alla igår . Det kommer gå fint . 
Hur många människor är det i det här rummet ? 
Om vi tar direkt perception som underlag för diskussion , som i Gibsons modell , skulle jag säga att jag uppfattar två personer , förutom mig själv . 
Så ... svaret borde vara tre . 
Försök igen . 
Hur många människor är det i det här rummet ? 
Hej . 
Allt bra ? 
Du såg inte pigg ut igår . 
Jag mår bra . Jag ville bara inte festa . 
Det är nog stress . 
Jag blir också glad när allt är över och vi kan fortsätta där vi slutade . 
Vårt sista år i frihet . Inte bara sitta och plugga . Vad är det för mening ? 
Lydia ? 
Vad sa du ? 
Efter det här kan vi leva som vanligt i ett helt år . 
Vad ? 
Är förändring alltid dåligt ? 
Det beror på förändringen . 
- Hur gick intervjun i dag ? 
- Dåligt , tror jag . 
Jag var bakis . 
Visste du att fresior symboliserar tillit ? 
Alltså , jag ... 
Jag tänkte att om jag lämnade Keshav ifred , skulle han få tid att komma till klarhet . 
Men han anpassar sig bara efter sina föräldrars åsikter . 
Han uppvaktar Camille ... och är inte sann mot sin verklighet . 
Och ... Jag borde inte ha släppt taget om honom . 
Det borde jag fan inte . 
Du hade kanske inget val . 
Det har man alltid . 
Man kan kämpa eller ge upp . 
Men varför är folk så rädda för att vara det de är ? 
Jag sätter mig längst bak och sover lite . 
- Ville du sitta här ? - Det är lugnt . 
Välkomna till studenternas frågestund . 
Jag lurade i mina klasskamrater att det fanns snacks och dricka här . 
Nu är de hungriga och känner sig lurade . 
Förhoppningsvis svarar de ändå på era frågor . 
Fråga på . 
Hur mastiga är kurserna här ? 
- Hinner man ha ett privatliv ? 
- Nila ? 
Det är mer intensivt än andra universitet . 
Det är sant , men oroa dig inte , man hinner ändå ha ett liv . 
Fler frågor ? 
Har man mycket kontakt med andra colleges här , eller är det separat ? 
Måste jag säga adjö till min bästis ? 
De är vanligtvis ganska åtskilda . 
Nån som har valt Balliol , till exempel , har inte så mycket att göra med nån som studerar vid St Hildas . 
Nej , Balliol är ju elit-colleget . 
Det är vad nån från Balliol skulle säga . 
Tack . Några fler frågor ? 
Vad är ditt betyg ? 
- Ursäkta ? 
- Jag undrar bara om du har kompetens att förbereda oss för detta . 
Vissa har riktiga frågor . 
Låt dem prata istället för att slösa tid på dina inkompetenta kommentarer . 
Har du problem ? 
Det är läskigt att du låter som han plötsligt . 
- Vem ? 
- Din far . 
- Ni kanske ... - Håll käften , din pajas . 
- Låt honom vara . - Förstör jag er dejt ? 
Varför är du här ? 
Du vill till Balliol , men låtsas inte att det var ditt beslut . 
- Vad ? 
- Det är din strategi . 
Du trycker ner och stöter bort alla , så att ingen märker att du bara är en fegis som går i ledband för att inte behöva stå för nåt . 
Ruby ! 
Du har ignorerat mig på sistone . 
Fortsätt gärna med det . 
Du har rätt . 
Jag går i pappas ledband , jag ljuger och döljer mina känslor . Men jag gör det för din skull . 
- Vad menar du ? 
- Glöm det . 
Prata med mig . Sluta prata i gåtor . Du gör mig galen ! 
Du gör mig galen ! 
Vet du vad du gör mot mig just nu ? 
Hur tror det känns för mig att höra din röst ? 
Du kan inte bara dumpa mig och skämma ut mig inför alla , och sen låtsas att jag missförstår . 
Jag kan inte ... 
Jag är ledsen , okej ? 
Vad gör du här då ? 
Varför pratar du med mig ? 
För att jag ... För att ... 
Du vet inte , för du vet inte vad du vill . 
Du vet ingenting ! 
Jag vet vad jag vill . 
Du kämpar inte för det . 
Ingen bryr sig om vad jag vill . 
Jo , jag . 
Det har jag alltid gjort . 
Du trodde väl inte på riktigt att nån som jag var intresserad av nån som du . 
Ruby ? Vad är det ? 
Jag är ledsen . Varför ? 
Vad är det ? 
Mina föräldrar märkte att du fick mig att förändras . 
Pappa såg dig som ett hot . 
Han hade rätt . 
Han svor på att han skulle förstöra ditt liv . 
Och jag kan inte skydda dig . 
Du förtjänar nån som kan skydda dig och en snäll svärfar . Det kan jag inte ge . 
Det enda jag kan erbjuda är en massa jobbiga problem . 
Varför sa du inget ? 
Du får inte bestämma åt mig . 
Han ville skada dig . 
Jag är inte rädd . 
Hur gör du ? 
Du vet inte hur han är . 
Jag vill inte ... 
Jag kan inte ... 
James . 
Sluta nu . 
Inga fler lögner . 
Jag lovar . 
Vad gör du ? 
Det par gör när de litar på varann . 
- Par ? 
- Du är inte min toy boy . 
Hur kan nån ha en så hög IQ och använda ord som " toy boy " ? 
Passar det att retas nu ? 
Jag är vad du vill . Pojkvän , toy boy , vad som helst . 
- Vad som helst ? 
- Allting . 
- Är detta killen som sabbar vattensängar ? 
- Det var inte en vattensäng . 
Jag stannar här . 
- Jag åker aldrig hem . - Du ville ju inte till Oxford . 
Jag sa inget om det här rummet . 
Vi stannar här . 
I morgon fortsätter världen gå runt . 
Du har lika många chanser som alla andra . 
Du måste använda dem . 
När jag är vilsen eller olycklig gör jag listor . 
Det motiverar mig och rensar tankarna . 
Gör du min lista ? 
Vad ska stå överst ? 
Jag gillar sport , musik ... 
Och stark asiatisk mat . 
Jag vill äta gatumat i Bangkok . 
- Friterade gräshoppor och så ? 
- Precis . 
Okej . 
Mer läsning ... 
Dessa är inte livsmål . 
Drömmar är viktiga . 
Jag mår bra när jag ritar . 
Önska dig nåt ! 
Du glömde det viktigaste . 
Miss Bell . 
Säg mig , varför Oxford ? 
Har ni hört om elefanten och stolpen ? 
En metafor för självbegränsande tankar . 
Att de flesta människor är kapabla till mer än de tror . 
Men jag börjar inse att jag har tjudrat mig vid min framtid . Och därför har många stunder i nuet inte fått den uppmärksamhet de förtjänar . 
James Beaufort ? 
James Beaufort , Balliol ? 
Nu vet jag att det är uppehållen vi gör på vägen som egentligen är livet . 
Livet här och nu . 
Och ibland kan dessa stunder rita nya spännande framtidsvisioner i sanden . 
Det här är Cordelia Beaufort . 
Lämna ett meddelande efter tonen . 
Hej , mamma . Jag hoppas att du mår bra . 
Jag har nåt att berätta . 
Oroa dig inte , det är ... goda nyheter . 
Jag älskar dig . 
Vi ses senare . 
Vi inser att vi inte fruktar framtiden längre . För det är nuet som avgör om våra drömmar ska bli sanna och om vi ska bli de vi alltid har velat bli . 
Det krävs mod för att tänka bortom nuet . 
Men ibland är det nån annans blick som kastar nytt ljus över vår framtid . 
För första gången kände jag att jag var framme . 
Hallå . Jag är hemma . 
Jag vill inte snabbspola framåt eller bakåt . Jag vill vara här , nu . 
Mr Beaufort väntar på er . 
Sätt er ner . 
Sätt dig , sa jag . 
Er mamma har fått en stroke . 
- Var är ... - Hur ... 
Cordelia är död . 
Vi åkte till sjukhuset , de kunde inte göra nåt . 
Och du ringde inte oss ? 
Cordelia var så stolt över er . Jag ville inte störa intervjuerna . 
Som jag sa är det vår första prioritet att hålla investerarna nöjda . 
Aktierna får inte gå ner . 
Ja , för satan , jag vet . 
Utkastet måste iväg . - Snarast . - James , nej . 
Ja för fan , Gordon , jag vet . 
n utses efter att pressmeddelandet gått ut . 
James , nej ! 
Sluta ! 
Rör mig inte ! 
Du satt i bilen och sa ingenting . 
Förlåt , James . 
Alla människor förtjänar en värld av möjligheter . 
Att drömma sina egna drömmar , att vara sig själva , att älska vem de vill . 
Jag ser min framtid tydligare än nånsin . 
Äntligen är alla pusselbitar på plats . 
Alla dörrar är öppna . Nu är det bara att gå genom dem . 
