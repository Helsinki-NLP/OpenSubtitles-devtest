- Sasà , han är skallig ! 
- Nej ! 
Han hade krulligt hår senast någon såg honom . 
Wonderboy ! Jag har bevis att han finns ! 
Munaciello har alltid funnits . 
Det är folket som har glömt att stan är full av magi , 
Vi har bara några dagar kvar tillsammans . 
Vi flyttar till Brescia imorgon . 
Inuti den här statyetten finns en skattkarta . 
Eftersom du inte gav mig statyetten , får du inte mina lägenheter ! 
Hyresvärden vill ha statyetten ! 
Hon kommer inte att ge efter för några krav från oss . 
Då gör jag det själv . Jag går in vid Gaiola . 
- Aniello , vad gör du ? - Aniello ! 
Aniello hoppade från klippan för vår skull . Vi måste rädda honom . 
Gaiola ... Neapels mest hemsökta plats . 
- Teresa ! - Teresa ! 
Du är Wonderboy ! Där är han ! 
Han har försvunnit ! 
Hör ni ? Såg ni Wonderboy ? 
Man ser ingenting här nere . 
Vi måste härifrån innan vi blir förkylda . 
Utan att hitta Wonderboy ? 
Vadå ? Skulle han rädda oss om vi hittar honom ? 
Ta det lugnt ! 
Vi ska träffa Clemente . Han skulle hjälpa oss ut . 
Vi måste bara ta reda på vart vi ska . 
Var är ungarna ? 
Så , du vill alltså bråka med mig ? 
Du vill lägga beslag på statyetten och lägenheterna . 
Vad snackar du om ? 
Det där bryr jag mig inte om . 
- Jag är här av en annan anledning . 
- Ingen bråkar med Capuozzo . 
Nu ska du ta dig ner och hitta statyetten . 
Du är verkligen galen ! 
Omöjligt . 
Vill du att jag ska slå mig fördärvad ? 
Föredrar du att dö så här ? 
- Är alla okej ? 
- Ja , men det är kallt . 
Du har en undervattensficklampa ! 
Jag kan inte ta mig ner utan redskap . 
- Se efter själv . Det är för djupt . 
- Så hur tar man sig ner ? 
- Rep och karbinhakar , grottutrustning . 
- Grottutrustning ... 
Okej . 
Ta den där ! 
Ta den . 
Ta den ! 
Titta där ! 
Är det vägen ut ? 
Vi ser efter . Kom igen ! 
Upp med dig , Aniello . 
Ge mig lampan . 
Vänta på mig ! 
Vi måste hitta Clemente vid mötesplatsen . 
Han väntar på oss ! 
Vilken väg ska vi ta ? 
Vi ser efter var den här tunneln tar slut . 
En genial plan . 
Vi har inget annat val . 
Kom nu . 
Oscar , titta här . 
Det här är Sasàs . 
Barnen har varit här . 
Är du säker på det här , Antò ? 
Ska vi gå in här själva ? 
Donna Angè , väggarna har rasat in ! 
Vi sitter fast ! 
Chihuà , var är du ? 
Donna Angè ! Jag hör dig inte ! 
- Vad händer ? 
- Han har stängt till ingången . 
Var är du , din idiot ? 
Jag tror inte det är sant . 
Kära nån , allt har rasat ihop . 
Sasà ? Var är du ? 
Ta dig ut ! 
- Maltè , sätt fart ! - Kom igen ! Vad gör vi nu ? 
Var är du ? 
Oscar , låt det vara . Vi kommer inte in här . 
Vad gör vi nu ? 
Vi berättar för alla föräldrarna och letar reda på en karta över gångarna . 
- Hjälp ! - Hjälp ! 
Vad händer ? 
Det är min pappa . 
Håll dig still , Dò ! - Kom ! Han kommer att hitta oss . - Ropa på honom . 
- Vad säger du ? 
- Vi måste härifrån ! Vi är vilse ! Nej , vi måste hitta Wonderboy och statyetten . 
Vi ville rädda dig . 
Har Chihuahua kommit hit för att rädda mig ? 
Hörni , vi måste röra på oss . 
Nu går vi . 
Seså , Rafè . Vi måste samarbeta . Kom nu . 
Långsamt , Enzo ! 
- Långsamt ! 
- Vad ser du ? 
- Ingenting . Det finns inget här . 
- Titta noga . 
- Vänta ! 
- Vad ? 
Jag ser något , men det är långt borta . 
- Det kan vara statyetten . 
- Ta den ! 
Det går inte ! 
All blod rusar mot mitt huvud . 
Dra upp mig ! 
Jag tar den från en annan ingång . 
Jag har kartor över Neapels underjordiska gångar i min husbil . 
Du sa att det här var enda vägen in ! 
Låt mig hämta andan . 
Hallå där ! 
Kom igen nu , killar . 
Brescia väntar på oss . 
Sätt igång nu . Det är dags att vakna . Vad är det med er idag ? 
Herregud . Var är de ? 
Snorungar . 
Var är ni ? 
Raffaele ! 
Gennà ! 
Var är de ? 
Nedrans snorungar ! 
Vad står på , Francesca ? 
Tvillingarna är försvunna . Alla är borta , Sasà och Teresa med . 
- De tog sig ner i underjorden . 
- De låg inte i sina sängar . 
De håller på med sina påhitt som vanligt . 
Hyresvärden är involverad också . 
Alla letar efter samma statyett . 
Är hyresvärden involverad ? 
Jag ska prata med henne . 
Vi ska till Brescia . 
- Lugna dig . 
- Francè , vad säger du ? 
Hon har aldrig hjälpt oss , och hon lär inte börja nu . 
Vi frågar Samantha . 
Hon kanske vet nåt . 
Hallå ! Samà ! 
Samantha ! Kom ut ! 
- Vad är det ? 
- Vad är Aniello och Chihuahua ? 
- De har gått härifrån . 
- När då ? 
Ingen aning . Jag har inte sett dem sen igår . Igår ? 
Var har de sovit ? 
Francè , det är inget ovanligt . 
Ibland är de borta i tre dagar . 
Vi är en modern , fri familj utan regler . 
Javisst . Men just nu kan de vara i fara . 
Barnen har varit nere i underjorden hela natten . 
- " I underjorden " ? 
- Neapels underjordiska gångar . 
De håller på med sina påhitt om stadslegender och gamla historier . 
Men de har inte kommit hem än . 
Hör du mig ? 
Fråga hyresvärden . Jag vet att hon vet något . 
Du är hennes frisör . - Ni är vänner . 
- Är du galen ? 
Jag stör inte henne för fyra ungars skull . 
Fem . 
Din unge är med dem . Har du glömt honom ? 
Hon är förbannad . 
Det har jag förstått . 
- Donna Angè . 
- Chihuà ! 
Klamra dig inte fast i mig ! 
Du drar ner mig ! Vad tror du att jag är ? En livboj ? 
Jag tror att vi är i en vattencistern . 
Och killen som stal statyetten ? Var är han ? 
Jag kan inte hitta honom . 
Han är nog död ! 
Och snart drunknar vi också ! 
Pitone ! 
Åk till Gaiola och hämta hit de där tre idioterna . 
Skynda på ! 
Varför är ni så värdelösa allihop ? 
Ni har blivit lurade av en kille i huvtröja ! 
Vem är han egentligen ? Spindelmannen ? 
Välkommen hem . 
- Har han sugkoppar på händerna ? 
- Gör han volter i luften ? 
Osynlighetsförmåga ? 
Hur kan han försvinna i tomma intet ? 
Jag sa ju det . Wonderboy kan allt . 
- Okej . Vad har du sett honom göra ? 
- Han klättrade som Tarzan och räddade mig . 
Såg ni inte hur han försvann i vattnet ? 
- Han kan ha drunknat . 
- Kom igen . 
Varför sa du så ? 
Vad är det för ljud ? 
Det låter som musik . 
Det låter som skräckfilmsmusik . 
Jag tänker inte gå dit . 
Vi går den här vägen . 
- Vart tar du vägen ensam ? 
- Var tysta ! 
Jag känner igen melodin . 
Terè , vi går härifrån . Vi ska gå upp , inte nerför . 
Det är beckmörkt ditåt , men där finns det ljus och musik . 
Vad ska du göra med lägenheterna ? 
Du kunde bett om vad som helst , men du valde hyreslängan . 
Och de är råtthål , värre än min husbil . 
Varför frågar du om det ? 
Jag är bara nyfiken . 
Nu förstår jag varför alla kallar dig för snåljåp . 
Är jag en snåljåp ? 
Jag föddes i de där hyreslängorna . Jag växte upp där , fram tills en dag ... då den där haggans föräldrar knackade på och sparkade ut oss . 
Nu vill jag få tillbaka vad som är mitt . Fattar du ? 
Jag ska rulla dem extra hårt , precis som du gillar . - Då varar de hela dagen . 
- Donna Angè . 
Hittade du dem ? 
Det har varit ett ras på Gaiola . 
Man kan varken ta sig in eller ut . Det är omöjligt . Vi måste hitta en annan väg att få ut dem . 
Tusan också ... 
Sluta med det där ! 
Säg åt Aspide att köra fram bilen . 
Vi ska åka till Andarnas slott . 
Vad är det som händer , donna Angè ? 
Handlar det där om min man ? 
- Samà , inte nu . - Ursäkta . 
Jag är orolig . Jag inte sett honom sen igår . 
Jag ska ta hand om det . Okej ? 
Låt mig göra klar din frisyr . Jag gör det själv . 
Nu räcker det . Jag ringer polisen . Vänta , Francè . 
Vad ska du säga till dem ? 
Okej . Jag går dit ensam . 
Hyresvärden är involverad . 
- Och Chihuahua också . 
- Har du hajat det nu ? 
Ni verkar lyda hennes order . 
- Du påstod att din familj var så fri . 
- Vi jobbar för henne . Det är annorlunda . 
Igår natt var hon på Gaiola och pratade med Clemente . 
Han som bor vid Andarnas slott . 
Oscar , berätta . 
De skulle åka dit nu , till Andarnas slott 
Ciro , hämta din van . 
Kom igen ! Vi måste hinna dit före dem . 
- Kolla upp det där . 
- Det här fixar jag . 
Vad gör du ? 
- Flytta bilen . Skynda på . - Ja , gärna . 
Jag ska på möte , men bilen vill inte starta . 
Vad är det nu ? 
Är du här , donna Angè ? 
Ursäkta mig . Det går inte en dag utan att den här rishögen bråkar . 
Idag är det bromsen som krånglar ... 
Vad nu ? 
Oj ! Vad är det här ? 
Hur kan det finnas ljus och musik här nere ? 
Mamma mia ... 
Den här melodin är så sorglig . 
Det är " Lu Cardillo " ... Det är en neapolitansk folksång . 
Mamma brukade sjunga den för mig . 
Du har rätt . Jag kände inte igen den först . 
Jag visste det ! 
Vi har upptäckt det här ! 
- Det är vi som är Wonderboys ! 
- Vad ? 
Det här är prinsen av Sanseveros hemliga laboratorium . 
Det här är en av hans största uppfinningar : " den eviga flamman " . 
Se här ... 
Inte ens vetenskapsmannen på tv kunde förklara hur den fungerar . 
Och här är speldosan . 
Det är som ett klockspel . 
Vad vackert det är . 
Varför vet du allt det här ? 
Jag läser mina läxor . 
Och prinsen av Sansevero var en stor man . 
I slutet av läroboken fanns det ett kapitel om alkemi som handlar om honom . 
Efter att han hade förlorat sin fru blev han galen . Han blev besatt av mysteriet om liv och död . 
Och så upptäckte han ett elixir som kunde väcka de döda till liv igen , " Aludel . " 
Det finns en formel , men ingen kommer ihåg var den finns . 
Okej , professorn . Vi fattar . 
Nu måste vi hitta vägen ut . 
Vad var det ? 
- Vad hände ? 
- Sasà , nej ! 
Nedrans ungar ! De är besatta i legenderna att de har dragit in den här stackaren . 
Ett knep som lärde jag mig i unga år . 
Så äckligt det är här . 
Prinsen av Sansevero skyddade sina uppfinningar och installerade fällor för tjuvar ! 
Milda makter ! 
San Severos anatomiska maskiner . Det här är inte sant ! 
- Wonderboy ! - Wonderboy ! 
Jag visste att du inte hade dött . 
Du är en superhjälte . 
Vad gjorde ni ? 
- Vad gör vi nu ? 
- Hur ska jag veta det ? 
Lugn ! Låt mig tänka efter . 
- Gennà. tänk snabbt ! - Ser ni vattnet där ? 
- Herregud ! 
- Hörni ! Snälla ... Hjälp ! 
- Vi måste hjälpa varandra ! Terè ... 
- Herregud ! 
- Aniè , kom ! Räck mig en hand ! - Hörni ! 
- Hjälp till ! - Hjälp ! - Vi sitter fast som i en råttfälla ! - Hjälp ! 
Tonì , du måste få ut oss härifrån . 
Är du ingen superhjälte ? 
Vad snackar du om ? 
Jag är här för statyetten . 
- Jag har inget med er att göra ! 
- Vad är grejen med statyetten ? 
Vad finns inuti ? Är det en diamant ? 
En skattkarta ? Vad ? 
Vem bryr sig om skatten ? 
Vi måste rädda oss själva . 
Gennà , hördu ... Prinsen satte ut fällor för att stoppa tjuvar ? 
Ja . Och det här är den bästa fällan . 
- Tjuvarna drunknar . 
- Det började när musiken slutade . 
Det måste vara nåt som en högtalare ... 
Eller en slags förstärkare ... 
Ser ni hålen i taket ? 
Vad menar du ? Går ljudet in där ? 
Just det ! Den uppfattar frekvenser och vibrationer . 
- När musiken slutar så triggas fällan . 
- Vänta ... 
Terè , du sa att du kan den här sången . 
Du måste sjunga den . 
Det är vår enda chans . 
Kom igen , Terè . 
- Terè , snälla . - Kom igen , Terè ! 
- Snälla , Terè ! - Snälla ! 
- Sjung , Terè . 
- Försök ! 
Sjung ! 
- Kom igen ! - Snälla ! 
- Vi ber dig . - Försök ! 
Men jag låter inte som en speldosa . 
Snälla . Det är vår enda chans . 
Snälla , jag ber dig . 
Oj ! 
Jag klarar inte mer . 
Kom , hörni ! Jag vet inte hur länge det håller sig öppet . 
Skynda er på ! Följ mig ! Kom ! 
- Skynda er på ! - Teresa . Hallå ... 
Kom igen . Kom . 
Teresa . Vi måste skynda oss . Kom nu ! 
Kom . Ner med dig . 
Kom igen , Terè ! 
Du har en fin sångröst . 
Det var sista gången du fick höra den . 
- Sätt fart ! 
- Okej . 
Nej . Nej ! 
Det har varit inbrott ! 
Nej . Den låg här ! 
Det var här jag lade den ! 
Enzo . De har stulit kartan . 
- Nu surnar jag till , Clemè ! - Nej , Enzo ! 
Lägg ner den där innan du skadar dig ! 
Antò , vänta ! 
Du är 18 , men vi andra är 40 . 
Snälla , berätta vart vi är på väg ! 
Antò , kan du förklara ? 
Ser ni korset ? 
Eftersom allt på Gaiola har rasat går vi in här istället . 
Och vad är det ? 
Det är en äldre ingång som har blockerats . 
Nu ligger den i villan där borta . 
- Vem äger den ? 
- Det Nino D ' Angelos villa ! 
Kom här . 
- Jag vill inte se dig igen . 
Okej ? - Vi är inte klara här ! 
Tack , Angè . 
Du räddade livet på mig . 
- Jag visste att du var en god ... 
- Var inte så dramatisk . 
Jag räddade dig för att jag behöver dig . 
Vad behöver du mig för ? 
Jag har några mannar som sitter fast under jord . 
Var är de ? 
Kom med mig . 
Var är vi nu ? 
Det är samma korsning som förut . 
Vattencisternen är därborta . 
Då så , hörni ... Nu säger jag hej då . Tack så mycket . 
" Hej då " och " tack " ? 
Vi räddade livet på dig och nu överger du oss ? 
Berätta vad det handlar om . Vi kan allt om Neapels gamla legender . 
Du vill ha statyetten för att hitta en gammal skatt , inte sant ? 
Nå , än sen ? 
Vi överlevde , eller hur ? Nu skiljs våra vägar åt . 
- Men vi måste ta samma väg . 
- Jaså ? 
- Låt mig vara ! 
- Nu tar jag hand om den här den här . 
- Maltè , ta honom . - Sätt fart . 
Donna Angè , hör du mig ? 
Donna Angè . Hör du mig ? 
- Chihuà ! 
- Vi har tagit tillbaka statyetten . 
Bra jobbat . 
Jag ska få ut er därifrån . 
Så vackert havet är idag . Hej . 
- Vadå ? Har du bråttom ? 
- Nej . 
Du har skyndat hit för att träffa mig ? 
Jag menar ... Det finns inget bra sätt att säga det här ... 
Nu blir jag nervös . Vad är det ? 
Jag är gravid . 
Du är gravid ? 
- Det är underbart , älskling ! 
- Ja , det är det . 
Vad nu ? 
Det är väl goda nyheter ? 
Ja , Alfrè . Det är bara ... 
- Vad ? 
- Mina föräldrar ... De kommer inte att acceptera dig . 
Det stämmer inte ! 
Jag tänker hitta skatten . Sen blir jag Neapels största filantrop . 
- Skatten . 
- Just det . 
Dina föräldrar blir stolta över mig och vi uppfostrar vårt barn tillsammans . 
Precis som i sagorna , okej ? 
Du är galen . 
Min baby . 
Donna Angè ... 
Ynglingen ... 
- Ska vi göra oss av med honom ? - Nej ! 
Jag vill träffa honom . 
Jag vill se honom i ögonen . 
Jag ska bevisa att Munaciello är en myt . 
