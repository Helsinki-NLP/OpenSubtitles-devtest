År 1946 Busan , Sydkorea Vi håller Busan under kontroll åt dig i valet . 
Nu räcker det . 
Vad läser du ? 
An Minchul Ledamoten An Yosubs äldste son 
Gillar du historieböcker ? 
Kang Seongmin , 16 år 
Varför läsa om kungar ? 
En kungason har bara två val . 
Han kan bli sin fars hund eller döda sin far och ta över tronen . 
Vad föredrar du ? 
Ingetdera . 
Hördu . 
Va ? 
Kom hit . 
Visa lite respekt för de äldre . 
Vill du inte bli kung måste du bli nåns hund . 
Din lilla snorunge . 
Vad sysslar du med ? 
Jag ber om ursäkt . 
Din son är modig . 
Han slog mig först . 
Din lilla ... 
Men han slog mig först . 
Vart ska du ? 
Jösses ! 
Vem är du ? 
Den dystra lilla jäveln . 
Är han din son ? 
Han är söt . 
Han är så deprimerande ! 
Så din mamma tog livet av sig här . 
Stirra inte på mig . 
Vad händer ? 
Din son dödade dig nästan , herr Kang . 
Fan ta dig . Kom hit . 
Kom hit , din odåga . 
Kom hit . 
Din lilla jävel ! 
När ska du ta ditt förnuft till fånga ? 
Du är som din mor ! 
Sineuialliansen står upp mot den makt som förtrycker vårt folk . 
- " Sineuialliansen står upp - " Sineuialliansen står upp - mot den makt - mot den makt - som förtrycker vårt folk . " - som förtrycker vårt folk . " 
Sineuialliansen kämpar mot orättvisa , och vårt våld är vår uppoffring . 
- " Sineuialliansen kämpar mot orättvisa , - " Sineuialliansen kämpar mot orättvisa - och vårt våld - och vårt våld - är vår uppoffring . " - är vår uppoffring . " 
Vårt första mål är Kang Ilsik . 
Kang Seongmin 
Cha Taemin , 25 år 
Uncle Samsik 
Uncle Samsik 
Hyckleri förklätt till en dröm 
Kim San går med i Demokratiska partiet som chef för ekonomiutskottet 
- Choo Intae ! - Choo Intae ! - Choo Intae ! - Choo Intae ! 
- Choo Intae ! 
- Tack , allihop ! 
- Tack ! 
- Choo Intae ! 
- Choo Intae ! - Choo Intae ! 
- Innovation är vårt hopp ! - Choo Intae . 
- Choo Intae ! - Choo Intae ! 
- Yeojin . 
- Choo Intae ! - Ursäkta mig . 
- Choo Intae ! - Dags för förändringar ! 
- Vad gör du här ? 
- Förlåt att jag dyker upp . Kan vi prata lite ? 
Inte nu . 
Vad vill du säga ? 
Jag tänker stötta herr Choo på nåt sätt . 
Att jag är demokrat förändrar inget . 
Ville du säga det ? 
Jag beundrar och stöttar herr Choo . 
Kan du gå ut dit och berätta att du är hans svärson ? 
Att du stöder Innovationspartiet ? 
Kan du lämna demokraterna ? 
Självklart . 
Yeojin . Du vet väl att jag älskar dig ? 
Jag har en dröm . 
Vad för dröm ? 
Jag vill förändra vårt land till det bättre . 
Det är ingen dröm . 
Det är hyckleri . 
Hyckleri förklätt till en dröm . 
- Choo Intae ! - Choo Intae ! - Choo Intae ! - Choo Intae ! 
Era jävlar ! Vad i helvete ? 
Yeojin ! 
Yeojin ! 
Snälla ... 
Yeojin ! 
Är du okej ? 
Hämta lite vatten . 
Varför var du där igen ? 
För att träffa Choo Yeojin ? 
Vårt avtal , då ? Jag måste väl förklara varför jag gick med i demokraterna ? 
Var inte löjlig . Titta på folkmassan ! 
Jag slutar . 
Jag har gett Yeojin så många löften . Jag måste hålla dem . 
Löftet du gav mig , då ? 
Är Choo Intae som din far och jag bara en farbror ? 
Varför är Choo Intae speciell ? Varför är han så bra ? 
Vad har han gjort ? 
Dessa nobla tänkare . 
De kunde inte ens ge sina barn mat under kriget ! 
Choo Yeojin vill inte vara politikerfru . 
Varför inser inte en smart man som du det ? 
Jag kan inte göra slut med henne så här . 
Varför inte ? 
Det är inte rätt . 
Vad skulle hon tro om mig ? 
Förutom pengar , makt och respekt , vill du vara snäll ? 
Du kan inte få allt . 
Jag slutar . 
Du är inte redo än . 
Jag kan ge dig pengar och makt , men jag kan inte även ge dig ära , kärlek och respekt . 
Jag bryr mig inte om det . 
Vill du höra min stora plan ? 
Åt helvete med den ! 
Hundra från liberalerna , 30 från demokraterna , tjugo som vinns över individuellt , plus 20 som kommer att nomineras i nästa val . 
Det är totalt 170 ledamöter , inklusive dig ! 
- Vi kan införa ett parlamentariskt system med den siffran . 
Oavsett vem som blir president , tar Cheongwooförbundet över nationalförsamlingen och utser premiärministern . Och det blir du . 
Aldrig att Liberala partiet stöttar mig ! 
Ja . De stöttar Kang Seongmin , inte dig . 
Han främjar systemet för att själv bli premiärminister . 
Vi får in dig i nationalförsamlingen inom tre år och utser dig istället för Kang Seongmin efter grundlagsreformen . 
Fokusera nu på ditt mål . Ditt nationella rekonstruktionsprojekt . 
Vill du bli premiärminister ? 
Svara mig . 
Ja . 
Lägg då all din uppmärksamhet på det du vill uppnå ! 
Jag vill göra det ! 
Jag vill genomföra nationella rekonstruktionsprojektet ! 
Jag gör slut med henne . 
Allt man vill ha i livet har ett pris . 
Håller du inte med ? 
Stanna här . 
Vänta . 
Är det inte säkrare med partimedlemmarna ? 
Ge mig bara en sekund . 
Jag går och kollar läget . 
Vad fan gör ni ? 
Du din ... 
Jag är er chef , idioter ! 
Din jävel . Hur dålig är du på ditt jobb ? 
Du är ingens chef längre . 
- Va ? 
- Slå mig , så är du dödens . 
Vad ska du göra ? 
Är du galen ? 
Slå mig om du kan . 
- Slå mig . - Hördu ! 
Gå . 
Låt mig göra det . 
Hallå där . 
Och vem är du ? 
- Flytta på dig , jävel . 
Ta dig samman . 
Jag löser det . Gå . 
Fan ! 
Herr Yoon . 
- Blev du skjuten ? 
- Ja . 
Du klarar dig , Haejun . 
Jongchul ! 
Haejun blev skjuten ! 
Jongchul ! 
Haejun , det är okej . 
Haejun ... 
Haejun . 
Hördu , Haejun ! 
Fan ! 
Haejun ! 
Fan ! 
Vänta utanför . 
Herrn ! 
Choo Intae blev skjuten . 
Va ? 
Vem blev skjuten ? 
Choo Intaes tillstånd är kritiskt . 
- Menar du allvar ? 
- Ja . 
Kritiskt tillstånd . 
Och Yoon Palbong ? 
Han dog på platsen . 
Jävla idioter . 
Ett vittne såg Cha Taemin från Sineuialliansen . 
Ursäkta ? 
Ja , vi undersöker det . 
Den avlidne är en gängmedlem vid namn Gu Haejun . 
Titta på det här . 
Fokusera ! 
Sail saltodlings 4:de chef Cha Taemin 
Ser du det här ? 
Jag gjorde det , eller hur ? 
Kom ut när du har skitit klart , idiot . 
Sluta skryta . 
Hej då , Haejun . 
- Efter dig . - Tack . 
An Yosub , vd för Segangs textilier , förlorade sin son i en explosion . 
Hans son var ledamot An Minchul , liberala partiets nya stjärna . 
Vem ligger bakom det ? 
Vem tjänade mest på hans död ? 
Kang Seongmin ? 
Cha Taemin från Sineuialliansen ? 
Fotot kan vara slutet för Kang Seongmin . 
Frågor om Sineuialliansen Terroristgruppen Sineuialliansen bakom Choo Intaes skjutning 
" Sineuialliansens våldsamma terrordåd är inte exklusiva för vänstern . " 
- " Vissa politiker ... " 
- Det är riktat mot mig . 
Ditt namn nämns inte . 
" En konflikt mellan politiker med affärsbakgrund . " 
De syftar helt klart på mig . 
Publicerades det med flit ? 
Bara Cha Taemin hade dessa bilder . 
" Explosionen i Busan kan vara relaterad till Sineui ... " 
Det räcker . 
Inrikesministeriet 
Vi organiserar grupper i varje departement och område och ändra lagen om lokalt självstyre . 
Så här går omröstningen till . 
Vi riggar 40 % av rösterna , och väljarna skriver in sig i grupper ... - Vad är det ? 
- Ta en titt . 
Som ni säkert vet från artikeln , är situationen allvarlig . 
Tror du att det är sant ? 
Har du sett bilden ? 
Det är väl Kang Seongmin ? 
Jag tror det . 
Varför skulle vi vara samlade om det inte var han ? 
Om ledamot Kang har varit inblandad i Sineuialliansen , behöver vi en plan B. 
I det här läget ? 
Det vore onödigt . 
Om Kang Seongmin får reda på det är vi illa ute . 
Oavsett om det är sant eller inte behöver vi en plan B. 
Enligt min åsikt borde vi göra en grundlig utredning först . 
Vi borde inte dra förhastade slutsatser och misstänka vår kollega . 
Jag gör några diskreta förfrågningar . 
Ja , presidenten . Ryktet verkar falskt . 
Artikeln var fabricerad . 
Ja , vi vidtar nödvändiga åtgärder . 
Ja . 
Partiet förbereder sig för att agera fortast möjligt . 
Är det sant ? 
Jag frågar dig , är det sant ? 
Det är inte sant . 
Jag blir förtalad . 
- Av vem ? - Jag undersöker det . 
Dödade Sineuialliansen ledamot An Minchul ? 
Jag vet inte . 
Det står så i artikeln . 
Det är bara ett antagande . 
Jag är säker på att An Yosub gör samma antagande . 
Utan Cheongwooförbundet är du värdelös . 
Jag ska döda den arroganta jäveln en dag . 
Nån kan höra dig . 
Hämta ledamot Pak Jiwook . 
Hej , herrn . 
Hej , herrn . 
Hej , herrn . 
Vad gör du här , herrn ? 
Har ni tagit Cha Taemin än ? 
Jeon Soyong Chef för nationella säkerhetsbyrån 
Han är svårfångad . 
Och Sineuialliansens övriga medlemmar ? 
De har varit inaktiva i över tio år . 
Du har väl en lista ? Ge hit . 
Varför skulle nationalförsamlingen ha det ? 
Ge mig den bara . 
Vi spårade dem för tio år sen , men fick släppa dem . 
- Varför ? 
- Ingen aning . 
Det var chefens order . 
Så mina män letar nog inte ens efter dem . 
Varför bry sig när de ändå släpps ? 
Samsik . 
Ja ? 
Vänta utanför , dr Hwang . 
Arbetade Kang Seongmin med Sineuialliansen ? 
Han växte upp med Cha Taemin i Busan . 
Vem dödade min son ? 
Cha Taemin eller Kang Seongmin ? 
Det vet jag inte . 
Hur mycket kampanjbidrag skickar vi denna månad ? 
Två miljoner hwan till nationella säkerhetsbyrån , tre miljoner hwan till inrikesministeriet , och fem miljoner hwan till Liberala partiet . 
Stoppa betalningarna . 
Okej , herrn . 
Hitta Cha Taemin och ta reda på vem som dödade min son . 
Ja , jag ska leta efter honom . 
Herr Cha . 
Herr Cha . 
Jag tog med lite mat . 
Och whisky . 
Och dessutom , här är lite pengar . Här är en båtbiljett från Busan till Shimonoseki om en vecka . Kolla tiden . 
Är Choo Intae ... död ? 
Det är inte säkert än . 
Choo Intae ... Jag ville inte döda honom . 
Oroa dig inte . 
Det är Yoon Palbongs fel . 
Göm dig bara . 
Kommer farbror Samsik ? 
Självklart . 
Vad sa An Yosub ? 
Han frågade vad som hände i Busan . 
Det är oroande . 
Ja , du . 
Var är Cha Taemin ? 
Varför frågar du det ? 
Kang Seongmin bad mig fråga dig . 
Han kom inte till vår träff . 
Var ska du träffa honom härnäst ? 
Varför skulle en ledamot vara så nyfiken ? 
Det är väl en vana från den japanska polisen . 
Du har rätt . 
Jag borde ha skjutit ihjäl dig när jag arbetade med den japanska polisen . 
Förlåt , herrn . 
När flyr Cha Taemin till Japan ? 
Nästa vecka . 
På ett fraktfartyg från Busan . 
Och biljetten ? 
Cha Taemin har den . 
Är han i Busan nu ? 
Jag vet inte . 
Den jäveln . 
Är du okej ? 
Ja . 
Detta är anledningen till att Yoon Palbong dödades , eller hur ? 
Kolla alla adresser . 
Skugga alla . 
Vad gör vi om Cha Taemin dyker upp ? 
Om ni känner er hotade , får ni döda honom . 
Var är han troligtvis ? 
Börja leta runt Kang Seongmin först . 
Har han verkligen nåt att göra med Cha Taemin ? 
Sluta ställa dumma frågor och gör som jag säger . Du vet bättre än så . 
Skulle vi träffa Taemin i fritidshuset ? - Ja . 
- Byt plats . 
Ledamot Kang , var du inblandad i Sineuialliansen ? 
Har du hört ryktet att du beordrade ett mord på ledamot An ? 
Verkar det vara jag på bilden ? 
Jag var inte säker själv . 
Förnekar du ryktena ? 
Förnekar du din inblandning i Sineuialliansen ? 
- Ledamot Kang ! 
- Har du inte pratat med media än ? 
Jo , men det funkade inte . 
Om jag är tyst tror alla att ryktena är sanna . 
Cheongwooförbundets kampanjbidrag har inte kommit än . 
Lite inte herr An på Kang Seongmin ? 
Det är absurt . 
Så varför har vi inte fått betalt än ? 
Kang Seongmin verkar ha förlorat hans tillit . 
Misstänker mitt eget parti mig nu ? 
Herrn . 
Varför beter du dig så här ? 
Ge det lite tid , så kommer pengarna . 
Hur vågar de säga så till mig ? 
Du borde träffa herr An innan ryktena sprider sig . 
Vad ska jag säga ? 
Be honom skona ditt liv eller nåt . 
Om Cheongwooförbundet inte skickar våra kampanjbidrag går inte lagen om lokalt självstyre igenom . 
Ilmos sjukhus 
Yoon Palbong hittad död 
Är herr Kim San inne ? 
San . 
Jag presenterade Yoon Palbong för Innovationspartiet . 
Hur kände du honom ? 
Vi arbetade tillsammans . 
Hans nyheter har oroat mig . 
USA:s militärdepå i Korea - Tack för ditt arbete . 
- Tack . 
Det ser bra ut . 
- Det ser bra ut . 
- Okej . 
- Tack . - Ingen orsak . Tack . 
- Njut av maten . 
Här . Tack . 
- Tack . 
- Det är inte mycket . 
Men det är för mycket . 
Att uppfostra fyra barn är inte billigt . 
Jag betalar mer sen . 
Behåll det . 
Tack , herrn . 
Tack . 
Jag ska träffa Oh Inwoo . 
Avsändaren är okänd . 
Finns det mer bevis på Kang Seongmins inblandning i Sineuialliansen ? 
Inte direkt , men ... Kang Seongmins far dog i en explosionsolycka . 
Sineuialliansen var kända för sina bomber . 
Titta vad jag hittade . 
Varför dödade Cha Taemin Yoon Palbong ? 
Enligt polisrapporten sköts Yoon Palbong först . 
Han var inte ute efter Choo . 
Hade Yoon Palbong nåt med Kang Seongmin att göra ? 
Jag tror det . 
Farbror Samsik . 
Oj , du skrämde mig . 
Vad gör du här ? 
Jag vill hämnas honom . 
Du vet vem som dödade Haejun , eller hur ? 
Känner du till Sineuialliansen ? 
Nej . 
De har mördat nyckelpersoner inom politiken på båda sidor . 
Det kvittar . 
De är extremt farliga . 
Det kvittar . 
Okej . 
Då är det nåt du måste göra . 
Jag gör vad som helst . 
Ilmos sjukhus 
Var snäll och gå . 
Följ din dröm . 
Att du sitter här är den värsta sortens hyckleri . 
Var snäll och gå . 
Gå bara . 
Har du hört nyheterna ? 
Ja , det är så synd . 
Är du redo nu ? 
Ja , herrn . 
Jag behöver ingen trevlig kille . 
Det här är en krigszon . 
Du behöver ett hjärta av sten . 
Jag tror att jag är härdad nog . 
Kan du besegra Kang Seongmin ? 
Det måste jag om jag vill överleva . 
Var Samsik var inblandad i mordet på Seodaemunligans Gu Haejun ? 
Jag vet inte . 
Mordet på Yoon Palbong från Dongdaemunligan , då ? 
Så vitt jag vet var det en olycka . 
Så en ligamedlem bara råkade gå med i Innovationspartiet ? 
Jag hörde att han såg upp till herr Choo . 
Samsik var inblandad i mordet på Choo Intae , eller hur ? 
Nej . 
Det var en olycka . 
Menar du att Choo Intaes död var en olycka ? 
Choo Intae , Yoon Palbong och Pak Jiwook . 
Allihop ? 
Jag vet inte om det var en olycka eller oundvikligt . 
Men återigen , det är väl så ödet är . 
Är det inte förrädaren Jang Doo-sik ? 
Jag försöker rädda dig . 
Det är inte ditt öde att dö än . 
Hur skulle du förändra mitt öde ? 
Samsik tror inte på ödet . 
Han bestämmer själv , och när hans plan går i stöpet kommer han på en ny . 
Han är fast besluten att forma världen . 
Det är hans natur . 
Har jag format den här världen ? 
Nej , världen formade mig . 
