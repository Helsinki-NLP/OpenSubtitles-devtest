Hej , sömntuta . 
Hungrig ? 
Gillar du inte pappas sång ? 
Visste du att Elvis hade en schimpans som husdjur ? 
Jag menar allvar . 
Han hette Scatter och brukade gå klädd i hawaiiskjorta och dricka whisky . 
Vänta i bilen . 
Pappa är strax tillbaka . 
Ska Anastasia flytta nu ? 
Ja , Kitty . 
Hon ska flytta till sitt nya hem . 
Får hon det bra där ? Självklart . 
Hon får det jättebra . 
Du måste vara " King " . 
Nåja , till affärerna . 
Gå inte för nära . 
Oj ! Henne var det fart i . 
Det gillar jag . 
Det är fart i dig . 
Eller hur , min skönhet ? 
Det här räcker inte . 
- Det är tio . 
- Vi sa 15 . 
Nej . Du sa 15 . 
Jag sa tio . 
Vad gör du ? 
Priset är 15 . 
Vet du egentligen vem jag är , herr King ? 
Du borde ta de tio . 
Men hej där , lilla damen . 
Är det din dotter ? 
Kitty , du skulle ju vänta i bilen . 
Förlåt , pappa . 
Nöj dig med tio . 
Kitty . 
Anastasia stannar hos oss ett tag till . 
Varje brottsfall är som en bok , med egna karaktärer och huvudhandling och bihandlingar . 
En utredning är som en samling av sidor ur en bok . 
En ledtråd här , en ledtråd där , som till slut måste jämkas samman för att skapa mening i det hela . 
Men man vet aldrig säkert om man har funnit alla sidorna . 
Eller om sidor ur en helt annan bok kan ha blandats ihop med dem . 
Ja , man kanske inte ens vet om boken handlar om en försvunnen prinsessa eller ett monster i skogen . 
Eller kanske båda ? 
Men man måste ändå skapa en trovärdig historia av det man har där alla delar och karaktärer i intrigen knyts ihop bra . 
En bra historia . 
Och det är lättare sagt än gjort . 
Okej . Var var vi ? 
Såg han dig ? 
Jag vet inte ! 
- Shit , shit , shit ! - Sluta säga shit ! 
Han är i källaren ! 
Han kommer att se dina tjejsaker ! 
Tjejsaker ? 
- Vad gjorde han där ? 
- Farmor ringde honom . 
Strömmen gick visst . 
Var det du som gjorde det ? 
Om jag inte använder hårtorken , blir håret stripigt . 
Herregud . Wanda ! Det är inte mitt jobb att se till att ingen märker att jag är inlåst i er källare . 
Okej , vi tar det lugnt , bara . 
Ingen panik . Bara ... 
Nej . 
Du måste svara . 
- Jag tänker inte svara . - Jo . Du måste tala med honom . 
Nej . 
Varför viskar vi ? 
Nej . 
Chris ? 
Tjena , kusin ! 
Läget , polarn ? 
Jag är i farmors källare . 
Du har visst dekorerat lite ? 
Ja , lite grann ... Du vet , bara för att göra det lite mysigare . 
Mysigare ? 
Är det nåt du inte berättar ? - Ljug inte för mig kusin . 
- Vad menar du ? Har du en flickvän ? 
Ja ! Just precis . Så är det . 
Du har alldeles rätt . Avslöjad ! 
Din Casanova där ! 
Okej , vem är hon ? 
Du vet ... En brud som jag har träffat . 
Du vet ? Inget allvarligt . 
Det är bara en tillfällig grej . 
Du fattar ? 
Ja , absolut , kusin . 
Häftigt . Det här måste firas . 
Jag trodde du skulle förbli oskuld . 
Ja , jättekul . Du skämtar . 
När får jag träffa den mystiska damen ? 
Snart . 
Snart , absolut . 
Är hon snygg ? 
Jaha ? Fega inte ur nu och var " bara vänner " . 
Du vet hur du är . 
Jag ringer dig imorgon . 
Här är Morgonnyheterna på Sundersheim FM - och vi har lite kusliga nyheter idag . 
I natt blev en lokal gymnastiklärare angripen av ett vilddjur ute i skogen , enligt uppgift ! 
Han är tydligen utom fara men fick några benbrott . Aj . Verkligen ? Ett vilddjur i Sundersheimskogen ? Eller hur ? 
Tror du att det kan vara ... - Nuppelwocken ! - ... Nuppelwocken ! 
Jag tänker då inte gå ut i skogen idag . 
Okej , nu ska vi lyssna på låt nummer tre på topplistan . 
Hej där , store man . 
Sovit gott ? 
Några pannkakor ? 
Gör du pannkakor ? 
Visst gör jag det . 
Får man inte göra pannkakor åt familjen ibland ? 
Hur var dataspelspartyt ? 
Du sov visst över hos Vinsons , sa mamma ? 
Vi borde ta bort buggarna därifrån . Jag visste inte att du kände dem så bra . 
Har ni buggat deras hus ? 
När då ? 
För en vecka sen , tror jag . 
God morgon . 
Oj , du gör frukost ! 
Hej , mästarn . 
Hur var Games World ? 
Bra . 
Toppen . 
Och hur mår Alex ? 
Du borde bjuda hit honom . 
Vi vill gärna träffa honom . 
Visst . Han är alltid välkommen . 
Hm . Pappa sa att ni satte kameror i deras hus ? 
- Varsågod , mon chéri . 
- Tack . 
Okej . Vad pågår ? 
Varför är ni så konstiga ? 
Har nåt hänt ? 
Är nån av er döende ? Nej , nej . 
Ingen är döende . 
Nej . Så ... Vi vet att vi på sista tiden har låtit saker bli lite ... Lite galna , kanske . Ja . 
Lite galna . 
- Det är okej . 
- Nej , det är inte okej . 
Vi saknar Wanda så mycket , men ... Men du är kvar här och vi är fortfarande dina föräldrar . 
Så vi lovar att försöka vara bättre . 
Mot dig och mot varandra . 
Vi vill bara att du ska veta att vi älskar dig mycket och alltid finns här för dig . 
Du kan lita på oss , okej ? 
Så , ska vi ge upp ? 
Nej . Nej . 
Vi ska aldrig ge upp . 
Men vi ska försöka låta bli att bli gripna , dödade eller angripna av vilda djur . 
Vi måste skydda familjen . 
Annars blir vi utskällda av Wanda . Ja . 
Ni vill ha en gruppkram , va ? 
Chris ? 
Du är vaken . Jag trodde du skulle sova hela dagen . 
Vad är det ? 
Inget . 
Jag visste inte var du var . 
Försökte du ... Nej . 
- Säkert ? 
- Vadå ? Nej ! 
Tänk efter . Efter allt som hänt , skulle jag bara sticka iväg ? 
Hoppas inte det . 
För du inser väl att om du rymmer är jag den siste du bör vara rädd för . 
När King inser att du är vid liv har vi båda en måltavla på ryggen . 
Och var tror du att de först letar efter dig ? 
Vill du att en sån som Lukas ska komma hem till dina föräldrar ? 
Har du kunnat sova ? 
Nej . 
Och du ? 
Jag är som en sengångare . Jag kan sova överallt . 
Har du sovit här inne hela tiden ? 
Det är inte så illa . 
Man vänjer sig . 
Jag hade glömt hur stort det är utomhus . 
Det är galet hur fort man vänjer sig vid saker , som hur en guldfisk aldrig blir större än sitt akvarium . 
Är den här ren ? 
Typ . 
Jag behöver borsta tänderna och håret . 
Det känns som att vara på en musikfestival . 
Fast utan musik . 
Och utan festival . 
Jag kom ihåg ett gammalt hus . 
Jag och polarna brukade gå dit som tonåringar när vi ville komma bort . 
Det är ett ödehus mitt ute i obygden . 
Vi borde kunna gömma oss där medan vi gör en plan . 
Nån stal den . 
Men ni anmälde det inte . - Nej . 
- Nån aning om vem som stal den ? 
Jag hann inte se så noga . 
En kort knubbig en och en lång mager en . 
Vad är buren till för ? 
Är den olaglig ? 
Vad gjorde ni igår bakom fru Wagners rododendronbuske ? 
- Det var väl uppenbart ? 
- Varför var ni där , herr Bartels ? 
Harald Hessel . Känner ni honom ? 
Nej . 
Han bor några hus från Wagners . 
Han verkar tro att nån spionerar på honom . 
Okänd för mig . 
Och hon ? 
Lenka Němková . Hon dog i en bilolycka i Tjeckien , 30 minuter från gränsen . 
Men 24 timmar tidigare var hon på Kapitän . 
Liksom ni . 
Samma dag som Wanda Klatt försvann . 
Dominik , saken är att du redan är villkorligt frigiven för innehav av ett stort antal olagliga ormar . 
Så om du skulle bli åtalad för ett annat brott , som att bajsa offentligt , sitter du i skiten . 
Obs vits . 
- Vad hände Nuppelwocken-kvällen ? 
- Jag vet inte . 
Var är Wanda Klatt ? 
Jag vet inte . Jag svär . 
Varför dödade du Lenka Němková ? 
Jag har aldrig dödat nån ! 
Jag kör åt King . Det är allt jag gör . 
- " King " ? - Ja . 
Förlåt . 
Här är listan du bad om . 
Alla återförsäljare i trakten som för kameror och övervakningsutrustning . 
Ursäkta . 
Jag säger inte ett ord till utan min advokat . 
Så om jag inte är anklagad för nåt , vill jag gå nu . 
Igår kväll blev en gymnastiklärare allvarligt skadad på en joggingtur , efter att ha angripits av vad han beskrev som ett " jättelikt odjur " . 
Jag är här med Hester Horn , - lokalhistoriker ... - Hej . 
... och organisatör av Nuppelwocken-vandringsturen . 
Fröken Horn , exakt vad är Nuppelwocken ? 
Den sågs faktiskt första gången redan år 717 , då Pippin den korte sägs ha träffat på besten under en ridtur i skogen . 
Monstret grep tag i Pippin , slängde in honom i buskarna och massakrerade hans häst tills bara benen fanns kvar . 
Man kan faktiskt se benen av hästen i mitt museum . Barn halva priset . 
En fascinerande historia . Och det finns säkert mer bakom . 
Ursäkta . Kan jag hjälpa er ? 
Överintendent Rauch . 
Har ni övervakningskameror ? 
Typ buggar , menar ni ? 
Verkligen lustigt . Ni är den andra som frågar efter buggar denna månad . 
Det måste vara nåt i vattnet . 
Vem mer frågade om dem ? 
En konstig familj . En grävling åt upp deras fåglar och maken ville göra en podd om det . 
Han kom tillbaka häromdagen med sonen . De köpte en sån där . 
Ingen dålig utrustning . 
Den ... Den är Oles . 
Ni vet , pojkar och prylar . 
Nå , fick ni reda på vad som hänt gamle Hessel ? 
Vi har inte funnit spår efter övervakningsteknologi hittills . 
Men om nån planterar ut buggar i stan , ska vi hitta dem . 
Vi har utrustning nu som kan kolla ett rum blixtsnabbt och hitta alla buggar . 
Verkligen ? 
Fascinerande . 
Men varför skulle nån vilja ta en sån risk ? 
Det är ju helt mot lagen . 
Jaha , på återseende . Japp . 
- Adjö . - Ja . 
Hon vet . 
Om de börjar söka efter buggar ... Ingen panik . 
Hon har inga bevis . I så fall vore vi gripna nu . 
Vi måste bara ta bort buggarna innan de hittas . 
Ta bort dem ? 
Hur ? 
Det var svårt nog att få dit dem . 
Vad ska vi säga ? " Hej , det är vi igen . 
Vi undrar om batterierna i er TV-fjärrkontroll behöver bytas ? " 
Om vi kunde hitta ett sätt att få ut alla ur sina hus några timmar ? Då kan vi ta alla i ett svep . 
Hur ska det gå till , Dedo ? 
Jag har en idé . 
Wanda Fest . 
Alla kommer att vara där . 
Alla hus är tomma . Vi kan gå in och hämta buggarna . 
Stå rakt , hakan högt , händerna ner . 
Starta musiken . 
Två , tre ... Ut med armarna . 
Och ner och till vänster . 
Inte höger , Nataly ! 
Och nästa position . 
Chassé . 
Selma , vännen , lätta steg , du låter som en elefant ! 
Och piruett . 
Och slutposition . 
- Carlotta . Dedo . 
Hej . - Vad tusan gör ni ? 
Vi väntade er inte idag . 
Ja , vi ville bara titta förbi och se hur det går . 
Tja , mycket är ogjort , men vi ska nog komma i mål . 
Jag insåg inte att det skulle bli så stort . 
Underskatta inte hur mycket Wandas försvinnande har påverkat stan . 
Vi undrade bara över tiden . 
Hur länge tror du att ni håller på ? 
Tja , om Jonas fick bestämma skulle vi hålla på hela dagen . 
Jag har redan sagt att han måste korta Sparkles från fem nummer till tre . 
Vi pratade om det och vill bara försäkra oss om att det inte känns framhastat . 
Ja , som vi ser det , - ju längre desto bättre . 
Okej . 
Då blir Jonas glad . 
Han var mycket besviken över att tvingas stryka sitt Kate Bush-solo . 
Det förstår jag . 
Vad gör ni ? 
Det är Beyoncé härnäst . Det där är fel kostymer ! - Jösses . 
- Ja . 
Jadå . 
Jag visste inte att så många människor var involverade . 
Ganska galet , va ? 
Wanda skulle ogilla det . 
Hon skulle slå ihjäl oss för att vi låtit det ske . 
" Ballonger ? 
Allvarligt ? " 
" Måtte de inte använda engångsbestick till buffén . " 
" Jag tycker att Jonas Vinson är skitjobbig . " 
Vi vet åtminstone att alla lär vara distraherade . 
En av oss måste ju vara här , det förstår du väl ? 
Efter allt de har ordnat för vår skull . 
Om Ole tar monitorerna och du tar buggarna , så måste jag klara av allt det här ensam . 
Det får inte hända . 
Vart ska vi ? 
Vi ska ordna med förstärkning . 
Tror du att det spökar här ? 
Kanske . 
Vad gör du ? 
Det brukade jämt vara ett fönster öppet här uppe . Jaha . 
Det var lättare när jag var 14 . 
Shit . 
Försiktigt . Jadå . 
Det gick bra ! 
Välkommen till min lya . 
Det är helgalet . 
Herregud . 
Funkar den än , tror du ? 
Vi tar reda på det . 
Undrar om det var de som bodde här . 
Ska vi dansa ? 
- Hej . 
- A-Alex . 
Tänker du inte be mig stiga in ? 
Visst . Absolut . 
- Kan jag ta din jacka ? 
- Tack . 
Vill du ha nåt att dricka ? 
Eller nåt att äta ? 
Vi har lasagne . 
- Nej tack . - Okej . 
Tänker du gå på tillställningen för din syster ? 
- Wanda Fest , menar du ? - Ja . 
Ja . 
Min familj går lätt till överdrift när det gäller såna saker . 
Jo , om igår kväll ... Ja , ingen fara . 
Jag ska inte säga nåt . 
Jag fattar . 
Vi var berusade . Det var ett misstag . 
Tycker du att det var ett misstag ? 
Jag menar , all alkohol och att jag spydde på den trevliga flickans skor . Det var väl inte idealiskt , precis . 
Och det andra ? 
Vadå ? 
Du menar , kyssandet och så ? 
Jag menar det är inget jag direkt ångrar . 
Ole , du måste ha bättre självförtroende . 
Jag menar , det är lite sött , men också irriterande . 
Jag visste inte att du var ... Jag trodde du var ... 
Jag är ingenting . Jag är ung . 
Jag behöver inga etiketter . 
Jag gillar dig , du gillar mig . 
Det är inte så komplicerat . 
Förklara för mig varför vi inte har bott här de sista tre månaderna ? 
Jag visste inte om det fanns el här . - Jag trodde att den var avstängd . 
- Nån betalar visst räkningen än . 
Voilà . 
- Skål . 
- Skål . 
- Vad är det ? 
- Jag hittar inte mobilen . 
Lugn , den är här nånstans . 
Lämnade du den i skåpbilen ? 
Hittade du den ? 
UPPRINGNINGAR LUKAS ( 19 ) Okej , ingen panik . 
Din lögnaktiga lilla skit . 
När jag hittar dig skär jag öronen av dig . 
Du är så gott som död , hör du det ? 
Du lär önska att du aldrig sett Wanda Klatt ... Okej , nu kan du få panik . 
Rüdiger , vi ville träffa dig för att ... Först och främst vill jag be om ursäkt för mitt beteende . 
Vill du ? 
Jag borde inte ha sagt det där till polisen , och du ska veta att du är en viktig del av vår familj , och att vi litar på dig och älskar dig . 
Jag älskar er också . 
Och förlåt att jag drev med din hästsvans och dina kläder och åkte hem till dig och klådde upp dig . 
- Du klådde inte upp mig precis . 
- Tja , det var rätt ... 
- Jag fick in några bra smällar . 
Ja , men sammantaget vill jag nog säga ... 
- Vi kan kalla det oavgjort . - Oavgjort ? 
- Jag fick in några bra snytingar ... - Okej ! 
Vi har stridit mer än nog . 
Så vi borde tala öppet om allting . 
Okej ? Det är en cirkel av tillit . - Okej ? 
- Cirkel av tillit . - Okej , jag börjar . - Ja . 
Jag miste jobbet men sa inget till Carlotta . Sen lånade jag pengar av dig och satte oss båda i en svår situation . 
För det vill jag be er båda om ursäkt . 
Min tur ? 
Okej . Jag köpte en tiger på mörka webben . 
En tigrinna , närmare bestämt , Klo-dia . 
Men hon kom aldrig och jag miste 26 000 euro . 
Hur kunde du köpa en tiger ? 
Du kunde inte ens hålla liv i kaktusen du fick på din födelsedag . 
Ska det inte vara en cirkel av tillit ? 
Det är sant . 
- Okej . 
Min tur nu ? 
- Precis . 
Okej . 
De senaste månaderna har vi i hemlighet försökt hitta Wanda , och olagligt spionerat på alla våra grannar med hjälp av övervakningskameror , också köpta på mörka webben . 
Va ? 
Va ? 
Han vet , Wanda ! 
Lukas vet ! 
Och om Lukas vet så vet King , och de kommer att leta efter oss ! 
Ta ett djupt andetag ! 
Låt oss tänka logiskt ett tag . 
Om du var Lukas och fick veta att jag lever , skulle du tala om det för nån ? 
Jag menar , King anlitade honom , inte dig . 
Om King är så farlig som du säger , lär inte Lukas ringa honom och säga : 
" Jo , du vet den där saken som jag lovade fixa ? 
Jag lyckades visst inte med det . " 
Ja . 
Du har rätt . 
- Han försöker fixa det själv först . - Ja . 
Jag borde gå och prata med honom . Kanske tar han reson . Övertala honom att följa med oss till polisen ? 
Chris , han är en psykopat ! 
Han är ändå min kusin . 
Är allt okej ? 
Jadå , allt är toppen . 
Skulle det vara problem ? 
Du måste vara skärpt . Du har jobb imorgon . 
Vi är en man kort . - Vem ? 
- Bartels . 
Vad har hänt ? 
Ursäkta , jag minns inte att jag inbjöd till frågor . 
Okej . 
Dit ska du åka . 
Imorgon . 
Jag återkommer om tiden . 
Häftigt . 
Så där . 
- Du är hemma . 
- Hej . 
Vi har inte ... Vi bara ... Hej , fru Klatt . 
- Hej . - Herr Klatt . 
Du kan säga Dedo . 
- Dedo . 
- Alex . 
Så trevligt att äntligen träffa dig ordentligt . 
Läget ? 
Jag är Rüdiger , Oles coola morbror . 
Alex . 
Okej . Vad har ni för er då ? 
Ingenting alls . 
Vi har prov imorgon . Ole hjälpte mig att plugga . 
Jag är inte så smart som han . 
Det känner jag igen . 
Var inte ledsen för det . 
I skolan finns alltid genier , och så såna som vi , visst ? 
Vi får leva på utseendet . 
Dags för mig att åka hem , - men trevligt att träffa er alla . - Ja . 
Vi ses snart , Alex . 
Vi ses snart . 
- Hej då , Alex . - Hej då . 
Jaha . 
Jag går till mitt rum . 
En trevlig grabb , verkar det . 
Ja , de kommer visst väldigt bra överens . 
De kysstes . 
Kysstes ? 
- Vänta , så Ole ... - Ja . 
Och alla de här är aktiva ? 
Vi har letat efter Wanda men tror att intendent Rauch vet om buggarna , så vi måste ta bort dem innan hon hittar dem . 
Planen är att göra det när alla är på Wanda Fest . 
Jag tar bort buggarna med hjälp av Ole , och här är operationscentret . Samtidigt håller Carlotta och du folk upptagna på Wanda Fest . 
Faktiskt en rätt bra plan . 
- Vi borde ge den ett kodnamn . 
- Det behövs nog inget kodnamn . 
Du behöver inte räcka upp handen . 
Så , Wanda Fest , är det uppträdanden och så ? 
Jag kanske ska sjunga en sång ? 
- Vilken bra idé . 
- Utmärkt idé . 
Fast jag vet inte om Vinsons redan har spikat programmet , så ... Jag tar med gitarren . 
Okej , Wanda ? 
Hör på . Om vi bara skulle fortsätta köra ? 
Vi kunde nog nå Grekland på tre dagar eller så . 
- Grekland ? - Ja . 
Chris , bli inte ledsen nu , men vi kommer inte att åka till Grekland ihop . 
Jag måste tillbaka till min familj . 
Wanda . 
Jag är så ledsen för att jag drog in dig i det här . 
Jag vet . 
Det är galet , jag menar ... De senaste tre månaderna har varit de mest påfrestande och galna i hela mitt liv . 
Men på vissa sätt har de också varit de bästa . 
Det är väl hemskt att säga så , men ... Nej . 
Jag vet ... Jag förstår egentligen vad du menar . 
Jag önskar förstås att inget av det här hade hänt . Men om inget av det här hade hänt hade jag inte fått tillbringa den här tiden med dig . 
Sjukt , va ? 
Du tänker säkert : " Oj , vad han snackar smörja . 
Först tillfångatar han mig och låser in mig i sin farmors källare , och nu säger han att han ... " 
Varför kysste du mig ? 
Först och främst för att få tyst på dig . 
Vad är det ? 
Alltså , om du fortfarande oroar dig , så gör inte det . 
Jag ger mitt medgivande . 
- Måste jag friskriva ... 
- Nej , nej . Nej . Det är inte det . 
Jag ... Bara , jag har aldrig ... 
Det är inget problem . 
Du lär dig fort . 
Hej , du har ringt Schellenberg . 
Lämna meddelande efter signalen . 
Det är en kungakrona . 
Jag trodde att hon ville spela en häftig drottning , men det är ingen drottningkrona utan en kungakrona . Den där King som Bartels nämnde . Han som styr över hela smugglingen av vilda djur . 
Lenka försökte avslöja honom . Därför lät han döda henne . 
Wanda måste ha sett nåt hon inte borde ha sett . 
Var det inte ditt jobb att hålla henne borta från oss ? 
Det är inte så enkelt när du skiter i buskarna hos folk och lämnar din skåpbil övergiven mitt i stan . 
Du nämnde King . 
Hon försökte sätta dit mig för den försvunna flickan . 
Jag hade inget med det att göra . 
Hälsa King att jag gjorde mitt och dumpade journalisten på andra sidan gränsen , men jag vägrar ta skulden för mordet . 
King uppskattar allt du har gjort för oss . 
Dominik . 
Alltså , Schelli , jag trodde ett tag att ... Jag har faktiskt en sak åt dig . 
Som ett tack . 
- Verkligen ? - Ja . 
Du kommer att älska den . 
- Vad är det ? 
- Vänta . 
Här . 
Öppna det . 
Öppna , bara . 
Sista beställningarna ! 
- En färdknäpp ? 
- Tack , hej då ! 
Hej då ! 
Wanda ? 
Wanda ? 
Wanda ! 
