Prins Zuko . Kejserliga gardet ska ta prinsen i förvar . 
- Va ? - Gardet ? 
- De är redan på väg . - Lugna dig , löjtnant Jee . 
Jag var på amiral Zhaos skepp och gick igenom ... bränsleförbrukningen . 
Löjtnant Dang och jag arbetade långt in på natten . 
Det kom ett bud till Dang . 
Drick upp , du . 
Jag hörde dem diskutera nya order . Från eldfursten själv . Han ska låta sitt personliga garde hämta hem prins Zuko för att åtala honom . För förräderi . 
- Förräderi ? 
- Är du säker ? Ja . Dang gav sina män order att möta gardet . 
I natt ? Då är han här när som helst . 
Det är Zhaos verk . 
Han har övertygat Ozai om att du vänt honom ryggen . 
Pohuai . Zhao har räknat ut att du befriade avataren . 
Prins Zuko , du måste genast ge dig av . 
Vänta med att starta motorerna . Undvik huvudleder . Res på natten . 
Far får inte tro att jag svikit honom . 
Nej , men nu måste du komma i säkerhet . Jag reder ut det med Ozai . 
Tack , löjtnant Jee . 
Ta hand om er , Ers Höghet . 
Jee anade inget . 
Det var lätt att få honom att svälja betet . 
Vad ska du säga till eldfursten ? 
Jag ska säga sanningen . 
Att prinsen satte sina egna behov framför sina landsmäns . 
Och att hans son var en förrädare . 
Spränggelatin . 
Prinsen ! 
Zuko . 
Nu måste jag framföra mina kondoleanser till general Iroh . 
Det kom säkert som en chock för honom . 
Zuko är ute på egen hand . Han var inte alls som jag trodde . 
Han verkade så ensam . 
Chockerande . 
Sokka , Aang fick kontakt med honom . Eller hur ? 
Jag insåg att Zuko och jag bär mycket på våra axlar . 
Jag har hela tiden varit orolig för att jag inte vet vad jag gör . 
Och det gör jag inte . 
Jag har inte lärt mig mer bändning och lär fortsätta göra bort mig , men jag har åtminstone mina vänner vid min sida . 
Precis . Team Avatar . 
Vad är det ? 
Titta ! 
Det norra vattenfolket ! 
Vi klarade det . Äntligen är vi framme ! 
De är här ! 
Välkommen till Agna Qel ' a , avataren . 
Det här är ... Vackert . 
Det är perfekt . 
Vi har väntat på er . 
Djuret är i goda händer . 
Vi tar honom till jakbuffelstallet . Det är en rymlig , uppvärmd grotta . 
- Se till att han får sjögräs . Massor . 
- Självklart . 
Välkomna . Jag är Arnook , det norra vattenfolkets hövding . Jag erbjuder er vår gästfrihet och vårt beskydd , i havsandens och månandens namn . 
Tack . Vi har verkligen sett fram emot det här . 
Det gläder oss att kunna välkomna en länge saknad bror och syster från södern . 
Det här är mäster Pakku , vår främsta vattenbändare . Och det här är min dotter , prinsessan Yue , stammens andliga ledare . 
Det är nåt jag måste berätta . Ni är i fara . 
Avatar Aang ... 
Det låter säkert vansinnigt , men i en syn jag såg blev ni attackerade . Vi vet . 
För några dagar sen fick våra spejare syn på en flotta från Eldnationen . 
Vi har haft ögonen på dem sedan dess . 
Vi är tacksamma för att du är här . 
Med avatarens krafter på vår sida ska vi ge dem en läxa de sent ska glömma . 
Medborgare , detta är en stor dag då vi välkomnar mäktiga allierade . Vi ska fira deras ankomst med en festmåltid . 
En festmåltid . Andarna har skyddat oss ... - Sluta stirra . - Va ? Jag kan inte . Det är nåt med henne . 
- Har vi träffat henne förut ? 
- Nej . Sluta nu innan de tror att du är störd . Mer än du faktiskt är . 
Jag ska inte vila förrän vi har hittat skurkarna ! 
Våra fiender får inte komma undan med ett sånt fräckt brott . 
Jag vet var vi ska börja leta . 
Jag vet vem som gjorde det här . 
Det var Ozai . 
Ozai har förlorat all sin mänsklighet . 
Han har blivit så besatt av att erövra världen , att han inte tål att nån kommer i vägen , inte ens hans eget kött och blod . Jag förstår . 
Mina sympatier . 
Då blir det jag ska säga härnäst en aning obekvämt . 
Eldfursten har gett mig den äran att leda en stor armada med order att erövra norr . 
Avataren är på väg dit , till vattenbändarnas sista stora fäste , så jag ska inta det . 
Förlåt mig , amiral , men du var inte den första tilltänkta för ett så viktigt uppdrag . 
Jag medger att jag har liten erfarenhet av strid . 
Men det betyder samtidigt att jag inte har nederlag bakom mig . 
Till skillnad från dig . 
Det räcker . Det räcker ! 
Eldfursten tycker att din prestation är undermålig . 
- Men jag vann ! 
- Du borde ha gjort slut på honom tidigare . 
Du får genomgå en ny prövning imorgon . 
- Du förstår väl att han leker med dig ? 
- Han kastade ett stenblock mot mig . 
- Din far vet redan att du är bäst . 
- Han vill inte visa det för dig . 
Låt honom tömma sina fängelser och bussa alla sina bändare på mig . 
Jag ska bränna dem alla tills han erkänner sanningen . 
Vilken sanning ? 
Att jag är den utvalda . 
Gå och prata med henne . 
Och säga vadå ? " Hej . 
Sokka , det södra vattenfolket . " 
Det är bara en tjej . 
Hon är prinsessa och andlig ledare . Hon sover på en tron och livnär sig på dagg och solsken . 
Lägg av ! 
Stuvade havsplommon . Min favorit . 
Är det gott ? Hur smakar det ? 
Som ... Som hemma . 
Katara ? Tack för att du hjälpte mig att ta mig hit . 
Det hade jag aldrig velat missa . 
Jag fick ju se världen tack vare dig . 
Jaha , smakar maten bra ? 
Den är utsökt . 
Du sa att du är helt självlärd . Ja , jag har kommit en bit på väg , men har mycket kvar att lära . 
Jag ville träffa andra bändare , särskilt vördade mästare som dig . 
Det måste ha varit svårt att vara avskuren från andra bändare . 
Eldnationens anfall berövade dig mycket . Liksom oss alla . 
Det värsta var att jag inte kunde göra nåt åt det . 
Det viktiga är att du överlevde . 
Det är det vi gör . Vatten är förändringens element . 
Vi vattenbändare har alltid anpassat oss efter livets flöden . 
Sök upp Yagoda imorgon bitti . 
Hon är en av våra bästa instruktörer och kan hjälpa dig . 
Tack , mäster Pakku . 
Vad sägs om hjortron ? 
Här har du . 
Tack ! 
Hjälp mig att äta upp det här . 
Kom igen . Det är gott . 
Vad tycker du ? 
Jättegott . 
Som barn gömde jag mig här när pappa hade möten med byns äldste . 
Han ville visa mig hur allt fungerar , eftersom det en dag blir mitt ansvar . 
Inte så värst kul . 
Jag gömde mig här med tanterna och fixade efterrätt . 
Du är bara en tjej . 
Tvivlade du på det ? 
Nej , jag tänkte bara att du är prinsessa och säkert ... - Högfärdig ? - Ja . Nej , menar jag . 
Jag trodde det , men du är vanlig . 
Eller inte vanlig , för det låter dumt . Jag borde sluta prata nu . 
Jag förstår . Där ute framstår jag som ... Men det är det alla förväntar sig . 
Missförstå mig inte . Jag står gärna i folkets tjänst , men ibland måste jag gå undan och ... Fixa efterrätt ? 
Jag fattar . 
Där hemma var det min plikt att skydda byn . 
Jag tog det på allvar . 
På för stort allvar , enligt Katara , men grejen var ... Det var ditt ansvar . 
Ja . Och om jag inte hade gjort det vet man inte vad som hade hänt . 
Det var ett löfte till min pappa , och det tänkte jag hålla . 
Men det hade varit skönt att slippa oroa sig ibland . Ibland vill man bara vara ... En pojke ? 
Hur känner jag dig ? 
Prinsessan Yue . 
De är redo för välsignelsen . 
Tack , Hahn . 
Du behövde inte lämna festen . En av prästerna kunde ha kommit . 
Det var inget besvär . Jag lovar . 
Det här är vår ismur . Den har stått emot attacker i hundra år . 
Hövding Arnook , får jag tala med vår broder från söder ? - Några stridsråd . - Från mig ? Vill du fråga mig om strider ? 
Du har nåt som vi saknar . Erfarenhet . 
Berätta om Eldnationens rustningar . Är de gjorda av metall ? 
Det sägs att de har taggar på axlarna . 
Inte metall , utan läder . Och inga axeltaggar numera . 
Resten av plutonen borde få höra det här . Kan du prata med dem ? 
- Visst . 
Berätta , avatar Aang . Vilken taktik tycker du är den bästa för striden ? 
Får jag föreslå att du leder den offensiva fronten ? 
Du kan gå i spetsen för attacken ... Luftbändning är mest inriktat på försvar . 
Vi brukar undvika konflikter . 
Men du är inte bara luftbändare . Du är avataren . 
Det är den enda bändningen jag behärskar . 
Det var därför jag kom hit . Jag hoppades att nån kunde lära mig . 
Men vi har hört det berättas om att du har räddat byar . Du har besegrat Eldnationens plutoner och bekämpat monster . 
Hur lyckades du med det ? 
Mina vänner hjälpte mig . Vi samarbetar . 
Det hade varit klokt att fokusera på träningen under resan . 
Vi kan visst inte räkna med avataren . 
Vatten är liv . 
Vattnet låter livet blomstra . 
Och läka . 
Mäster Pakku sa att vi skulle få besök idag . 
Jag är tacksam . 
Jag visste inte att vattenläkning fortfarande användes . 
Ja . Det är en viktig del av vår kultur . 
Känn energin flöda genom kroppen . 
Koppla det flödet till energin inom dig . 
Läkning är inte bara en fysisk process . 
Det handlar om empati . 
Du måste förstå vad det innebär att känna smärta , och sen avlägsna den . 
- Du är en naturbegåvning . 
- Tack . Jag har fått lära mig saker snabbt . 
Vi har tvingats improvisera en del . Ett eldklot som närmar sig gör en fokuserad . 
Apropå det . När börjar vi med stridsträning ? 
Ursäkta ? 
Jag klarar grundformerna bra , men precisionen måste bli bättre . Och kraften . 
Kvinnor strider inte . 
Våra krafter läker . De tillfogar inte skada . 
- Jag vill inte bara göra det . 
- Läkning är en ädel och helig tradition . - Det högsta kallet av alla . - Nej , förlåt . Jag menade inte så . 
Men jag tror att mina färdigheter är bättre lämpade för strid , så om det går bra vill jag träna stridsteknik . 
Hos det norra vattenfolket får kvinnor inte delta i strid . 
" Får inte " ? 
Det är inte rätt . Men så är det . 
Uppfattat . 
Vilken bra grupp . 
Vi har lärt upp dem så gott vi kan , men ingen av dem vet vad som väntar . Ingen har upplevt en strid . 
De klarar det säkert , speciellt med dig som ledare . 
Jo ... Prinsessan Yue . Hon verkar toppen . 
Hon är hängiven , snäll och generös . 
Hon representerar våra högsta ideal . Hon är den bästa av oss . 
Du gillar henne . 
Prinsessan och jag var trolovade . 
Det arrangerades när vi var barn , men när hon blev 16 bröt hon förlovningen , vilket hon har all rätt att göra . 
Men hon angav inget skäl . 
Men hade du fullföljt det ? 
Tack för att du visar avatar Kuruk din vördnad . 
Jag vill göra mer än så . 
Jag hoppas att Kuruk kan hjälpa mig i striden . 
Är det ett problem ? 
Det var länge sen nån bad Kuruk om nåt . 
Minnet av honom har bleknat . 
Han var inte så engagerad i omvärlden som avatar . 
Han blev tydligen förtjust i Andevärlden och tillbringade den mesta tiden där . 
Det betydde tyvärr att han inte fanns här för att hjälpa oss med våra problem . 
Han skötte alltså inte sitt jobb som avatar . Han svek alla . 
Det är nog inte hela sanningen . 
Jag hoppas det , för jag behöver hjälp och han är den enda som kan förstå min situation . 
Hej , Aang . 
- Du har tagit dig norröver . 
- Ja , för det norra vattenfolket är i fara . 
Avatar Kyoshi visade mig en syn där Eldnationen hade ödelagt Agna Qel ' a . 
- Jag måste förhindra det . 
- Det kan du inte . 
Om hon visade dig ett ödelagt norr , så kommer det att bli så . 
Men vi vet inte hur striden slutar . 
Om Eldnationen går segrande ur den och om vattenbändarna överlever ... Det hänger helt på dig . 
- Jag är bara ett barn . 
- Nej , du är avataren . På Kyoshi-ön hjälpte avatar Kyoshi mig att släppa loss otroliga krafter . 
Avatartillståndet . 
Ja ! Det gav mig samma styrka som tusen bändare . Med den kraften kan jag rädda norr . 
Men för att få kontroll över den måste du bemästra de andra elementen . 
Men hon kunde ta kontrollen . 
Hon kunde kanalisera kraften genom min kropp . 
- Hon hade kontrollen . Du kan göra så . - Det går inte . 
- Jo . Kyoshi gjorde det . - Jag är inte hon . 
- Du kan ändå göra det ! - Nej ! 
Efter att jag blev avatar upptäckte jag att mörka krafter var nära att ta sig över från Andevärlden till vår värld . 
Jag måste stoppa dem och lade hela livet på att bekämpa dem . 
Mitt krig mot andarna skadade min kropp och fördärvade min själ . 
I det här skicket kan jag inte bemästra avatartillståndet bättre än du . 
Och trots alla mina uppoffringar kunde jag inte rädda den som betydde mest . 
En rovlysten ande ville hämnas på mig . 
Ummi , min älskade , fick betala priset . 
Anden stal hennes ansikte . 
- Koh . - Lyssna på mig , Aang . 
Avataren måste vandra ensam . Annars får de du älskar lida . 
Ursäkta . Jag letade efter Katara . 
Jag ska väl gå , då . 
Är nåt på tok ? 
Nej , jag är bara lite trött . 
Du måste väl få töcknet att klarna . 
- Jag visste det ! Det var du ! 
- Ja . - Du är räven ! - Ja . Men hur ? 
Ganska snart efter att jag föddes blev jag mycket sjuk , så min far bönade och bad andarna att rädda mitt liv , och ett mirakel inträffade . 
Månens ande besvarade hans böner och gav mig en del av sin essens och räddade mitt liv . 
Det var då mitt hår bytte färg . Är du en ande ? 
Delvis , men mest människa . 
Jag tillhör båda världar och har varit en bro mellan dem . 
Jag blev prästinna för att hjälpa andra att få kontakt med sin andlighet . 
Det betyder att jag kan besöka Andevärlden . I mina drömmar . 
- Går du dit för skojs skull ? 
- Skulle inte du göra det ? 
- Det är magiskt . 
- Jag skulle välja ett annat ord . 
- Gillade du det inte ? 
- Om jag gillade det ? 
Att nästan bli sargad av ett monster , få ansiktet uppätet eller återuppleva smärtsamma minnen ... Smärtsamma ? 
Det var inget . Strunt i det . 
Gör inte så . 
Förminska det inte . 
Det var nåt som hände när jag var liten . 
Jag hörde pappa säga att han var besviken på mig . Att jag inte dög som krigare . 
Han trodde inte på mig . 
Vet du vad jag minns om dig från Andevärlden ? 
Du var orolig för dina vänner . 
Ditt hjärta . 
Det är det som utmärker dig . Det gör dig till en krigare . 
Om din pappa såg dig nu skulle han nog hålla med . 
Jag måste fråga en sak . 
Varför avvisade du Hahn ? 
Hahn är underbar . 
Han är allt en tjej kan önska sig . Men han är inte pojken i mina drömmar . 
Mina vänner betyder allt för mig . Jag klarar mig inte utan dem . De hjälpte mig hit . De kan hjälpa mig att vinna striden . 
- Vi är Team Avatar . 
- Det finns inget sånt . 
Det finns bara en avatar . 
Sluta tänka på vad du behöver och börja tänka på deras bästa . 
Att vara avatar innebär att man axlar bördan . Ensam . 
En björn ! 
Det är faktiskt en fisk . Den har en fena . 
Hallå . Pratade du med Kuruk ? 
Kan han hjälpa dig ? 
Nej , det kan han inte . 
Jag får klara mig själv . 
- Katara , hur gick det med Yagoda ? 
- Bra , men jag har en fråga . Var ska jag vara under striden ? 
Kvinnor får inte delta i strid . Jag trodde du visste det . 
Nej . Då hade jag inte godtagit det . 
Det handlar inte om att godta . Det är bara så det är . - Det är dumt och fel . 
- Det är inget att diskutera . 
Jag har slagits mot eldbändare sen vi åkte . Har dina män gjort det ? 
- Det kvittar . - Varför ? Det handlar inte om dem , utan om dig . 
Kvinnor är inte starka nog . 
Du har inte tränat och förberett dig på att ge ditt liv för alla andra . 
Vi ska inte gå samma öde till mötes som det södra vattenfolket . 
Jag får inte strida . 
De har varit instängda bakom sin mur så länge att de har fastnat i tiden . 
Vi kanske borde prata med Yue . 
- Eller ... - Vi kanske borde lyssna på dem . 
Du kanske inte borde strida . 
Den här striden blir inte som de vi redan har varit med om . 
Jag vill inte förlora er två . 
- Du kommer inte att förlora oss . 
- Men blotta tanken kan bli ett hinder . Människorna här behöver avataren . 
Jag kan inte vara avataren om ni är där . 
Jag undrar vad de kallar mig när nyheten når huvudstaden . 
Jag gillar " Zhao Erövraren " . Det ska låta lite slagfärdigt . Amiral , om jag inte misstar mig planerar du ett frontalangrepp mot staden . 
Staden är omgiven av oöverstigliga hinder på tre sidor . Framsidan skyddas av en ismur . 
Vad får dig att tro att du kan lyckas när andra har misslyckats ? 
Jag har nåt som de andra saknade . 
Jag har ödet på min sida . 
Vår propaganda hävdar motsatsen , men vattenbändarna är varken svaga eller fega . 
Om man underskattar dem kan det få tragiska konsekvenser . 
Otänkbart . 
Flottan har utrustats med nya , dödligare vapen , och vad viktigare är har jag personligen vidtagit åtgärder för att säkra vår seger . Vad är det ? 
Det här ... Det är ödet . 
Han ska angripa fästet framifrån , som en brunstig tjur . 
Mer vill han inte avslöja . 
Jag har underskattat Zhao . Han är farlig . 
Jag förstod det när jag simmade från min brinnande båt . 
Vi är snart framme i norr . Har du en plan ? 
En plan ? 
Planen är att visa att det var rätt av far att ge mig uppdraget . Och att fånga avataren en gång för alla . Och att återta det som är mitt ! 
Ingen plan , alltså ? 
Jag jobbar på det . 
Zhaos djärvhet förvånar mig . Det trodde jag inte om honom . 
Det känns nästan som om han jobbar med nån annan . 
Nån mycket smartare . 
Välj en motståndare . 
- Du måste välja en ... - Nej . Jag är klar . - Azula , sluta fåna dig . - Det är inte jag som fånar mig . 
Det är sista chansen . Ta striden eller bli underkänd . 
Att du bara vågar ! 
Vill du testa mig ? 
Släpp loss mig då . 
Släpp ut mig i världen , så ska jag visa vad jag går för . 
Jag har lekt färdigt . 
Pakku är en idiot . 
Det kvittar vad andra tycker . Det kvittar om pappa trodde på mig som krigare . Jag kan ändå vara bra på nåt sätt . 
Grejen är att det är min sak att avgöra , precis som det är din sak att avgöra vem du är . 
Jag ska utmana Pakku på en duell . 
Jag vet . Han är en mästare . Han sopar säkert banan med mig , men det spelar ingen roll . 
Jag har hållit igen hela livet . Jag tänker inte låta nån stå i min väg nu . 
Katara . Minns du när du sa att vi måste följa med Aang ? Att vi måste hjälpa honom ? 
Du hade rätt . 
Om vi inte hade gjort det hade jag inte vetat att två ungdomar från söder kan mäta sig med alla . 
Eldbändare , jordbändare , andevarelser , till och med stiliga krigare från norr ... Om du försöker prata vett i mig , så går det dåligt . 
Va ? Vadå , prata vett ? 
Nej , jag försöker säga åt dig att ge honom spö . 
Vad händer ? 
- Jag tänker inte slåss mot dig . 
- Du är bara rädd för att ha fel . 
Snälla . Gå tillbaka till läkehyddorna med de andra kvinnorna . 
Okej . Vill du lära dig att slåss ? 
Studera detta . 
Har du fått nog ? 
Var det allt ? 
En sak ska du veta . Du är en skicklig vattenbändare . 
Men jag får ändå inte strida . 
Ingen har pressat mäster Pakku så ! 
Det var otroligt ! De där isskivorna ... Hur gjorde du ? 
Kan du visa mig ? 
Nu kan ingen påstå att du inte är stark nog . 
Nej , bara att jag förlorade . 
Gjorde du ? 
Du sa att vi inte kan strida för att du inte vill förlora oss , men det är mitt beslut att strida , inte Pakkus eller ditt . 
Precis . Tror du att vi kom ända hit för att överge dig ? 
Din dummer . 
- Jag vet inte om jag kan skydda er . 
- Det kan du inte . 
Och att oroa sig för vem som blir skadad ... Det är inte bara avataren som gör det . 
Så är det att ingå i en familj . 
Kuruk , Roku , Kyoshi ... Alla sa att jag måste göra det på egen hand . 
Avataren måste axla bördan ensam . 
Det är historia . Bara en person kan berätta om framtiden . Den som ska skriva legenden om Aang . 
Hon menar dig . Det fattar du , va ? 
Eldnationen är här . 
Dags att ta strid . 
