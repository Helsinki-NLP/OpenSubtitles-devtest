Han måste ha lagt den där . Vem annars ? 
Tror du att Rusty la den där ? 
Vem annars vore desperat nog ? 
Mår du bra , Tommy ? 
Hon är rädd , jag bär upp henne på övervåningen . 
Hej , vad har hänt ? 
Va ? 
Har den testats i labbet ? Ja . Varken dna eller fingeravtryck . Troligen skrubbad . 
Hur vet vi att det här verkligen är Carolyns eldgaffel ? 
Det vet vi inte . Men kanske ni . 
- Dra åt helvete . - Och vi har det här . 
Det bevisar ingenting . 
Det bevisar att nån försöker skrämma mig eller sätta dit mig . 
Att nån föraktar mig . Det visar på nåns desperation . 
Vill du ta med den som bevismaterial ? Hur ? 
Det finns ingen förvarskedja , den är inte friande bevisning . Den kan bara beskrivas som " en eldgaffel " , inte " eldgaffeln " . 
Hushållerskan , då ? Kan hon identifiera den ? 
Vi tog hit henne . Den ser likadan ut , säger hon , från samma uppsättning , men mer kan hon inte säga . 
Och ditt hem har gåtts igenom ? Ja . Varken dna eller fingeravtryck . Lämnade inga spår . 
Inbrott ? 
Nej , jag lämnar sidodörren öppen . Jag har en katt . 
Ibland när jag jobbar sent kommer grannen över och ser till henne . 
- Ja . - Okej . Låt mig tänka . 
Jag är beredd att ogiltigförklara rättegången . Igen . 
Vad säger ni ? 
Åklagarsidan fortsätter gärna . Men vi anser att juryn bör underrättas om situationen . 
Vi kan låta dem veta att den inte ska ses som bevismaterial . 
Caldwell , då ? 
Varför skulle Caldwell vilja sätta dit Tommy ? 
- Ni gjorde honom förbannad ... - För att flytta fokus från dig . 
Domaren , jag behöver en stund med min klient . Tack . - Tack , domaren . - Det är en dum fråga . Visst . Förhörde ni honom ? Jag vill bara veta . 
Rusty , lugna ner dig . Rusty ... Det är så ... Lugna ner dig . 
Vi vill inte ha med det här , inte ens att det nämns . 
Med eller utan instruktioner . 
Men det kan så tvivel . 
Varför skulle Tommy ta fram det här om han inte talar sanning ? 
Att eldgaffeln är i hans förvar stärker ju inte hans fall . 
Och en lapp med texten : " Dra åt helvete " ? Det känns planterat . 
När sa du senast som åklagare : " Titta , jag hittade mordvapnet i mitt kök . " 
Instämmer . Det försvagar fallet . Och om vi vill bibehålla Liam Reynolds som en möjlig gärningsman , - talar detta mot det narrativet . - Okej , så nu vill du bibehålla Liam Reynolds ? - Inget motiv att sätta dit Tommy . - Vi borde fråga Caldwell . 
- Varför skulle han sätta dit Molto ? - Jag ... Vem vet ? Vem bryr sig ? 
Det handlar inte om sanningen , utan om att etablera rimligt tvivel . 
Lyssna på mig . Om juryn tror att eldgaffeln planterades , vilket de lär tro , misstänker de inte Caldwell , utan dig . 
Så de tänker inte nämna den alls ? 
Det är ju inte godtagbart som bevis , vilket kanske är lika bra . 
Det vore graverande för mig , för jag har motiv . 
Tänk om det läcks till media ? 
Jag menar , om det är till åklagarsidans fördel , varför skulle inte Tommy läcka det ? 
Om det kommer ut ogiltigförklaras rättegången , vilket han nog inte vill . Han tror att han ska vinna . Och de vet inte ens om det är mordvapnet , enligt dig . 
Det är det . Det saknas en flisa i handtaget . Jag kände igen den . 
- Berättade du det för dem ? - Nej . 
Jag använde den en gång där för att göra upp eld . 
Tur att inte mina fingeravtryck fanns på den . 
Vad är det ? 
Kan du ta ut den här ? 
Jag kommer strax . Jadå . 
Om en person äter och dör inom cirka 20 minuter finns det mesta av maten osmält i magen . 
En del går till tolvfingertarmen , inkörsporten till de nedre inälvorna . 
Fanns det mat i Carolyn Polhemus mage - när hon dog ? - Nej . 
Hur lång tid tar det för en människomage att tömmas ? 
Vätskor och liknande lämnar magen ganska snabbt , på mindre än två timmar . Proteiner och fetter cirka , 2,5 timmar . Ris och bönor , cirka tre timmar . 
Kvittot , stämplat kl 20 : 27 , visar kyckling kung pao och krabba rangoon som levererades till ms Polhemus hem kl 20 : 55 . 
- Ja . - Och när hon dog - var hennes mage helt tom ? - Ja . 
Ändå fann dr Kumagai att hon dog omkring kl 22 : 00 . Han har fel . Jag menar att hon dog mellan kl 01 : 00 och 03 : 00 . 
Hur kan han ta så fel ? 
Vet inte . För att hennes mage skulle vara tom måste hon ha dött minst fyra timmar efter att hon åt . 
Hon kanske aldrig åt maten ? 
Hon beställde den , den anlände . 
Kan du utesluta att nån annan kom ungefär vid den tiden och dödade henne innan hon hann äta ? 
Det fanns en halvfull behållare med kinamat i köket , så ... Fann du några spår av kinamat i hennes tolvfingertarm ? 
Det fanns spår av mat i tolvfingertarmen . 
Kan det ha varit hennes lunch ? Jag antar att allt är möjligt . 
Kan du fastslå med medicinsk säkerhet att offret åt kinamat ? 
Tack . 
Bara så att allt är klart , du jobbar enbart som expertvittne för försvaret ? 
Du har avgett en rapport med en åsikt , och därefter beslutar försvarssidan om de ska anlita dig eller ej , och om din åsikt inte gynnar försvarssidan , - anlitas du inte ? 
- Jag är professionell . Ett professionellt försvarsvittne som bara får betalt om dina åsikter gynnar försvaret och din åsikt idag gäller tiden för döden baserat på maginnehållet , där du antar att offret åt kinamat kl 22 : 00 . 
Har jag fattat rätt ? 
Okej . Låt oss anta att vi idag lyckades få juryn att tro eller åtminstone överväga att Carolyn mördades vid midnatt eller nån gång därefter . 
Vi måste bevisa att du var hemma då . Kan vi det ? 
Ja . Jag kan gå i god för honom . 
Vi kan inte kalla henne . Varför inte ? 
För att du är partisk och för att du ger dem tillfälle att utmåla din man i ett negativt ljus . 
" Stämmer det , mrs Sabich , att du inte visste att han låg med offret ? " 
" Stämmer det inte , mrs Sabich , att han fortsatte affären trots att han sa att den var slut ? " 
" Stämmer det inte att han inte berättade för er var han befann sig mordkvällen ? Att han gjorde henne gravid ? " " Hade ni en öppen relation , mrs Sabich ? " 
" Vet han allt om er ? " 
" Vi har alla våra hemligheter . 
Känner han till Clifton , den vänskaplige kvartersbartendern ? " 
Vad i helvete ? 
Har ni skuggat mig ? 
Ibland anlitar vi privatdetektiver enligt teorin att sanningen hjälper oss . 
Ibland gör den det . 
Vi avstår . Vi har rimligt tvivel . Varför ta risken ? 
Jag håller nog med . 
Jag tar slutanförandet . Åh nej . 
Nej . Det motsätter jag mig . 
- Det är mitt liv . Jag bestämmer . 
- Rusty , du har noll trovärdighet hos juryn . 
Varför skulle de tro ett enda ord du säger ? Alltså , jösses . I Maine , min hemstat , om en matar grisarna så måste nån annan mota dem . Jösses . Jag tar avslutningsanförandet . Om juryn tvivlar på mig , gör det inget . Om mina advokater tvivlar på mig , är det en helt annan sak . Eller om min bäste vän tvivlar på mig . 
Du borde kliva av . 
Det är inte möjligt . 
Klart att det är möjligt . Om han vägrar att följa dina råd ... 
Domare Lyttle låter mig inte kliva av nu . Det skulle anses påverka juryns utslag . 
Han är inte frisk . 
Frisk eller inte , oskyldig eller inte , han kommer att vara redo . 
Raring , den här rättegången har nästan dödat dig redan . 
Efter det här går jag i pension . Jag lovar . Jag ska ta promenader , klippa gräset , dricka iste med dig , bli rena Thornton Wilder och älska det alldagliga men vi är långt därifrån just nu . 
Det saknas bevis , vare sig fysiska , rättstekniska eller från vittnen . 
Nico Della Guardia ... Vi har också Liam Reynolds Caldwell , andra outredda jag från början offer . Så , jag gjorde det . 
Det är precis det ... Aldrig under mina 15 år som åklagare i vår fina stad har jag nånsin ogiltigförklarad rättegång , känslor för offret . 
Det hade jag med . Jag älskade henne mycket . 
Jag saknar henne mycket , och jag vill veta vem mördaren är , liksom många andra . Och jag förstår ... Hej . Hej . 
Jag övar på mitt slutanförande . 
Jag ser det . 
Behöver du hjälp ? 
Jag läste astronomi i skolan , så jag ser nog om nåt är från en annan planet . 
Et tu , min dotter ? 
Han blev lite galen mot slutet , du vet . 
Du vet , bli förrådd av sina vänner ... 
Sånt påverkar en . 
Pappa , allvarligt ? Slutanförandet ? 
Sa din mamma åt dig att komma in hit ? 
Jag är min bästa chans , Jay . 
Det här är mitt jobb . 
Jag klarar det . 
Bara några saker . 
Börja inte säga att Tommy är den verkliga mördaren eller Liam Reynolds , eller ex-maken . 
Hör du mig ? Rusty ? 
Ja , jag hör dig . 
Okej . 
Då är det försvarssidans tur . 
Mitt namn är Rusty Sabich , som ni redan vet . 
Jag är den anklagade . 
Anklagad för mord . 
Smärtan att tvingas säga det här i rättssalen inför min fru och mina barn ... 
Vad bevismaterialet klargör är att jag svek min familj , de människor jag älskar mest . 
Jag kan aldrig gottgöra den vånda jag har vållat min fru , och mina barn får troligen aldrig tillbaka respekten för mig . 
Men vad bevisen inte visar är att jag dödade Carolyn Polhemus , för det gjorde jag inte . 
Jag hade en affär med Carolyn , som jag hemlighöll . 
Jag gjorde henne gravid , vilket jag inte visste förrän efter hennes död . 
Och jag var där den kvällen som andra kvällar , men det är allt bevismaterialet kan visa , eller har visat . 
Det fanns inga ögonvittnen , det fanns inget blod eller rättstekniska bevis på mig eller på mina kläder , i min bil , i mitt hem . 
Mina fingeravtryck finns i hennes hem , för jag var där den kvällen som andra kvällar , men det är allt som kunnat bevisas . 
Tommy Molto stod här vid rättegångens början och sa att han hade känslor för offret . 
Det hade jag också . 
Jag höll av henne mycket . 
Jag älskade henne mycket . 
Och jag saknar henne mycket . 
Och jag , liksom många andra , vill veta vem som gjorde detta . Jag vill ta fast den skyldige . 
Liksom polisen och distriktsåklagaren , Tommy Molto . Han vill det så hett , att trots att han inte är säker , nöjer han sig med det näst bästa , nämligen mig . 
Och jag är som klippt och skuren . Omständigheterna pekar på mig . 
Det medger jag . Men inte bara på mig . 
Det fanns andra som var fixerade vid Carolyn . 
Vi har Michael Caldwell , offrets son , som också var där den kvällen . Och som var väldigt , väldigt arg på sin mor . Och som hade tillgång till Bunny Davis akt . 
Inte heller hans far , Dalton Caldwell , som också var väldigt arg på offret och som möjligen hade tillgång till Bunny Davis akt . 
Bevisar något av detta att Michael Caldwell eller Dalton Caldwell dödade Carolyn Polhemus ? 
Självklart inte , men nog måste man undra . 
Jag är åtalad . Jag är partisk . 
Men jag kan säga att under mina 15 år som åklagare i denna fina stad , har jag nånsin väckt åtal mot nån utan att bevisbördan är helt uppfylld , vilket är exakt vad åklagarsidan har gjort . 
De har åtalat mig för ett brott , men de har absolut inget som bevisar min skuld . 
Det finns inga fysiska , rättstekniska bevis , eller fällande vittnesmål . Det finns inget mordvapen . 
Det finns andra möjliga misstänkta som inte utretts . 
Och lägg till det Liam Reynolds , som öppet hotade offret . 
Och tiden för offrets död är oklar . Så det finns massor av rimligt tvivel . 
Så frågan bör ställas varför vi alls är här ? 
I fall med hög profil är det åklagarens plikt , som förresten är politiker , att tillfredsställa allmänheten . 
De måste ställa nån till ansvar . De måste hitta en ansvarig . Vem som helst . Och i det här fallet passar jag bäst . 
Jag är Tommy Moltos bästa chans . Han har velat fälla mig ända från början . 
Hans ogillande , hans förakt , har varit fullt synligt . 
Han har en agenda . 
Det här fallet . Det handlar inte om Tommy Molto eller om mig , eller ens om Carolyn , åtminstone inte ifråga om rättvisan , utan om er . Ni svor en ed att uppfylla en plikt , att för fällande dom får det inte finnas rimligt tvivel . 
Jag accepterar ert förakt . 
Jag förtjänar det . 
Och ... Som make ... Som far ... 
Men jag dödade inte Carolyn Polhemus , och därför finns inga bevis för min skuld . 
Jag är inte hedervärd . Men det ironiska är att jag hoppas att ni är det . 
Tack . 
Svaranden talade om sin kärlek till offret , men vad som har kommit fram under rättegången , och det mr Sabich medgav , inte bara var kärlek . Det var en fixering . 
Han sa att han ville hitta den skyldige . 
Men som vice chefsåklagare hade han alla möjligheter till det . Han ledde faktiskt utredningen . 
Jag kan tala om att de första 48 timmarna efter ett mord är avgörande för brottets lösning . Vad gjorde han under denna kritiska tid ? Han undanhöll information , han obstruerade , han befallde chefsutredaren att bara dela bevisning med honom själv . Och särskilt inte med mig . 
Han underlät att avslöja att han hade en sexuell relation med offret , att han var upprörd efter ett traumatiskt uppbrott , att han var i hennes hus mordkvällen . 
Han teg om allt detta . 
Så gör inte en oskyldig man , särskilt inte en vars plikt det är att gripa hennes mördare . 
Han ljög . Han dolde . Han försökte muta och utpressa andra att avge falska bekännelser . 
Han angrep vår rättsläkare fysiskt och slog ett potentiellt vittne . Så gör inte en oskyldig eller en som är mot våld , vilket svaranden påstår sig vara . 
Hans egen goda vän , Eugenia Milk , sa att han inte var sig själv dagarna innan mordet , utan gick helt upp i Carolyn . 
Han skickade 30 sms dagen hon mördades , inklusive detta : " Vem fan tror du att du är ? " " Vem fan tror du att du är ? " 
Han var där , han blev sedd där , hans DNA och fingeravtryck finns där , och ändå säger han på fullt allvar , med sin charmiga framtoning ... Han säger : " Det finns inga riktiga bevis . " 
Jaså inte ? 
Svaranden är en mycket skicklig lögnare . 
Och en mördare . 
Se vad som gjordes med henne . 
Dagen han åkte dit , dagen han sms:ade henne , dagen hon avvisade honom , och kvällen han sågs senast med henne , se vad som gjordes . 
Men han ställer sig och säger : " Det kan ha varit Liam Reynolds , det kan ha varit hennes ex-man . " 
Han antydde visst också att det kan ha varit jag . Det kan ha varit jag . Jaha . 
Det där är helt vanlig desperation . 
Det är normalt . Vad som inte är normalt är att han anklagar hennes son mitt i allt detta . 
Det är diaboliskt . Det är sociopatiskt . 
Hör på , svaranden hade som åklagare möjlighet att gripa personen som mördade Carolyn Polhemus . 
Men vad gjorde han ? Han dolde . Han obstruerade . 
Varför ? 
För han visste att mördaren inte fanns där ute nånstans . 
Mördaren fanns precis här . 
Det finns ännu en chans att skipa rättvisa , och den faller på er . 
Okej ? 
Han har gjort mitt ... Vad kallade han det ? 
Mitt förakt ! 
Mitt förakt , mitt uppförande till en faktor i sammanhanget . 
Okej . Han ber er att se på mig . 
Se på mig . Ta en ordentlig titt . 
Men också ta en ordentlig titt på den mannen . 
Det här är det värsta . Väntan . Eller näst värst . Att förlora vore nog ännu värre . 
Inte vet jag . 
Precis . Du är för bra för att förlora . 
Jag antar det . 
Allvarligt , hur ska vi tolka det ? Väntan ? 
Ju längre juryn överväger , desto mer gynnar det försvaret . 
Lika bra att vi går hem . 
Juryn kan dröja ett bra tag . 
Och jag oroar mig verkligen , för katten . 
- Ska det vara roligt ? - Det var ett skämt , Tommy . 
- Det är som att ... - Jag vet . ... vänta på att pannan ska koka . Vi går och tar en drink eller nåt . 
Jag tror att det var hans försäkring . Hela tiden . 
- Vadå ? - Eldgaffeln ? Okej ... Om han blir fälld , har han nåt att exploatera för en ny rättegång eller ... På nåt sätt . Jaha . Tror du att Rusty lämnade eldgaffeln i ditt hus ? 
Jösses , vad fan såg hon hos honom ? 
Får jag ställa en personlig fråga ? 
Hur mycket älskade du henne ? Allvarligt . 
Hör ni , domslutet . 
Jaha . 
Stå upp , mr Sabich . 
Vill rättsbiträdet läsa upp domslutet . Ja , fru ordförande . 
" Illinois högsta domstol , Cook County , i fallet åklagarmyndigheten i Illinois mot Rozat K. Sabich , fall nummer 6710098 , vi i juryn finner svaranden Rozat K. Sabich " " icke skyldig till mord " " i strid mot brottmålsparagraf 609.195 , ett grovt brott mot Carolyn Polhemus , en människa , enligt punkt ett i informationen . " 
Det känns overkligt . 
Det är över , va ? 
De kan inte överklaga eller begära ny rättegång ? 
Åklagarsidan överklagar inte . Det är över . 
Men ju förr de hör från mig , desto fortare sticker de . 
Jag är förstås nöjd med utslaget . 
Juridisk rättvisa skipades . Liksom moralisk rättvisa såtillvida att jag är oskyldig till det här brottet . 
Men rättvisa har inte skipats helt i det här fallet . Rättvisa har inte skipats för Carolyn Polhemus . 
Hennes mördare är ännu fri , och mordet är ännu olöst . 
Rättssystemet , särskilt åklagarämbetet , har svikit Carolyn Polhemus . 
Hon förtjänade bättre . Mycket bättre . Anledningen till att hon inte fick det var att de som anförtrotts att skipa rättvisa var motiverade av ärelystnad , och som jag misstänker känslor . 
Tommy Molto . Han hade skygglappar från dag ett . Han tappade målet ur sikte . Han hade redan bestämt sig , och distriktsåklagarämbetet misslyckades skändligen . 
De satte en vendetta före sanningen , och de svek framför andra Carolyn Polhemus . 
Tommy , du skötte dig utmärkt i rätten . 
Verkligen . 
Vårt fall byggde på indicier , och du gjorde ditt bästa . 
Han besegrade mig . 
Jag svek henne . 
Hennes död förblir ohämnad , för jag räckte inte till . Nej . Tommy , hör på . 
Du måste gå vidare . 
Det här är Chicago . 
Här finns en massa härligt avskyvärda skurkar att ge sig efter . 
Vi måste gå vidare och göra vårt jobb . 
Och själv behöver du släppa Rusty Sabich . 
Verkligen . 
Vi har jobb att göra . Låt oss sätta igång . 
Vi kan nog ta den där semestern nu . Du har visst packat . 
Det var dr Rushs råd om det skulle hända igen . 
Hända igen ? Ja . 
Om du nånsin mer skulle krossa den här familjen med ett impulsivt slag . 
Hända igen ? 
Jag visste egentligen från början , och sen visste jag inte . 
Men sen visste jag säkert . 
Rusty , jag vet inte vad du pratar om . 
Jag kunde bara tänka : " Det är mitt fel . Skulden är min . " Och jag gjorde vad jag måste för att skydda min familj , skydda dig . Vilket jag gjorde . 
Det som inte stämde var att du verkade så totalt normal nästa dag . 
Bara missnöjd . Jag visste inte att du kunde döda nån och vara så lugn . 
Tror du att jag dödade Carolyn ? 
Nej , det var nån annan , men nån i din kropp , liksom det nog var nån annan i min kropp som band henne . 
Menar du att du band henne ? 
För att skydda dig . 
Va ? 
Jag återvände samma kväll . 
Vad ... Först tänkte jag ringa larmcentralen , ifall hon möjligen var vid liv än , fast hon uppenbarligen inte ... var det . 
Sen slog det mig . Bara en person kunde ha gjort detta . 
Så jag ringde inte larmcentralen , för att skydda denna person , så att inga misstankar skulle riktas mot henne . 
Men allt det där med Liam Reynolds ? 
Falska bekännelser är lätta att framtvinga . Vi gör det ofta . 
Vi ... Jag erbjöd honom sänkt straff , vilket brukar räcka . 
Det var värt att pröva . 
- Rusty , du är sjuk . - Men sen började jag tänka : " Herregud , jag måste ta fel . " 
Men så berättade Jaden om dissociation , hur man kan bli avskild från jaget och stänga in en handling i ett fack , skilt från en själv . 
Då började jag inse att det var detta som hade hänt . 
Du tappade besinningen mot Carolyn , och nästa dag var det som om nån annan hade begått handlingen . 
Du är galen . 
Och du har fel ! 
Jag har inte fel . 
Efter din flört med bartendern spårade jag din bil . 
Va ? 
Jag vet att det var du som åkte till Tommy Moltos hus med eldgaffeln . 
För att hjälpa mig , antar jag , men du åkte dit . 
Nej , det gjorde hon inte . 
Det var jag . 
Va ? 
Jag ... Jag trodde att du skulle bli dömd efter ditt vittnesmål . 
Det var det enda jag kunde komma på . 
Vänta . Vad ... Jag körde dit i mammas bil . 
Va ? 
Jag la eldgaffeln i hans kök . 
Nej . Hur kunde du ha eldgaffeln ? 
Jag åkte dit för att konfrontera henne , och ... Hej . 
Vill du inte ha lite te ? Nej . 
... säga åt henne att lämna dig i fred . 
Lämna vår familj i fred . 
Det är inte jag , utan din pappa . 
Han vägrar lämna mig i fred . 
Det är inte sant . 
Du måste sluta ditt jobb och hålla dig borta från min familj för alltid . Håll dig borta . 
Jag ska hålla mig borta . Men hans liv och mitt kommer att vara lite sammanflätade . För jag är gravid med hans barn . 
Sen körde jag hem , och trodde att allt bara var en dröm . 
Men det var det inte . 
När ni åt frukost sa jag att jag inte mådde bra , och jag rengjorde bilen 
och grävde ner eldgaffeln . 
Okej , hör på mig . 
Vi ska aldrig prata om det här . 
Lyssna noga , Jay . 
Det här var nåt som kom ut ur dig som ett slags självförsvar . För att försvara den här familjen . 
Och det var jag som satte allt i rörelse . 
Jag bär skulden till det här . 
Vi ska överleva som familj . Okej ? 
Vi älskar varandra . 
Vi är en familj , och vi älskar varandra . 
