Det är bara jag , Kenny . Det är bara jag , Kenny . 
Major ? Överste Harding söker er . Ja . 
Allt väl , major ? 
Vi kommer alla att sakna major Cleven , sir . 
Väderrapport . 
Det tros klarna upp . Jaha , bra . 
Skjuts , major ? Nej , det behövs inte . 
Säkert , sir ? 
Bara lugn , Kenny . Jag känner inte av spriten . 
Vi ses imorgon . 
Bremen var det tuffaste uppdraget under hela kriget för mig . 
Den kraftigaste luftvärnselden jag nånsin hade upplevt . 
En granatskärva stor som en fotboll for genom planets nosparti och halshögg nästan mig och Douglass . och halshögg nästan mig och Douglass . 
Vänstervingen tog eld och vi miste all elkraft , men på nåt sätt fick Ev Blakely oss tillbaka till England . 
Jag såg också major Clevens plan ta en direktträff och störta . 
Från dagen jag anslöt mig till 100:e var Buck Cleven vår ledare . 
Vi såg honom som oövervinnlig . 
Om Gale Cleven inte klarade sig , vem kunde då göra det ? 
Kan vi hjälpa er ? 
Ja . Ni kan börja med att ge er iväg från vår förläggning . 
Och var är mitt skåp ? Va ? 
- Ursäkta , sir . De sa att ert plan ... - Men det gjorde det inte . 
Ta er utrustning och gå , mina herrar . 
Jag ordnar en ny barack . 
Ni har väl inte skickat hem mitt skåp redan ? 
Ni har väl inte skickat hem mitt skåp redan ? Nej , sir . Det är kvar i ordonnansens barack . 
Jag behöver en drink . 
Bra idé . 
Kom igen . 
Alltså , Dougie vad har du i ditt skåp som du är så orolig för ? 
Jag har tamejfan fler kondomer än jag kan räkna . Jag vill inte att min mamma ska räkna dem . 
Lugn , jag ska prata med henne . 
Titta , det är Blakelys besättning . 
Jösses , vi trodde att ni var döda . 
Fyra fallskärmar rapporterades från ert plan . 
Nån kan inte räkna . Det var ingen som hoppade . 
Via och Yevich är på sjukhus . 
Vi miste Saunders . 
Var landade ni ? 
Ett RAF-flygfält utanför Ludham . 
- En jäkla läskig buklandning . 
- Verkligen . Två motorer borta , hela flygkroppen full av hål . 
En mekaniker räknade . - Hur många var det , 1 200 ? - Tolvhundra . Stabilisatorn var paj . Landningshjulen gick inte att fälla ner . 
Landningshjulen gick inte att fälla ner . Men ingen fara , bromsarna funkade än . Tills vi landade . 
Rena undret att killen här , Everett Blakely , lyckades landa planet . 
Nej , undret var Croz bäring . En grad fel , så hade vi hamnat i vattnet . 
- Ren tur . - Du gör det för ofta för att det ska vara tur . 
Sen lyckades han styra oss rakt på det enda trädet inom synhåll , så ... Fullträff . En naturbegåvning . Det enda trädet i East Anglia , - och det träffar han . - Det största fältet ... - Harry Crosby ... - Rakt på . ... den bäste navigatören i 8:e flygflottiljen , där har ni honom . Vem är törstig ? Jag bjuder . Crank också . 
- Gör jag ? - Ja , det gör han . Kom . - Om du säger det så . - Härligt . 
Okej , kompis . - Bubbles ... hur mår du , kompis ? 
- Är det verkligen du , Croz ? 
Jösses , varför ringde du inte ? 
Det fanns ingen telefon på basen . 
- Men en lastbil som tur var . 
- Otroligt . 
Jag skrev till Jean . Du ... Ursäkta , vad gjorde du ? Jag skrev till din fru . Alla trodde att du ... - Du har väl inte skickat det ? - Nej , då . Tack och lov . 
Jag kom inte på nåt snällt att skriva , så ... Jag trodde faktiskt också att jag var död några gånger . 
Jag trodde faktiskt också att jag var död några gånger . Ja , men du klarade dig hem . 
Inte en dag för tidigt . De börjar göra förändringar i operationsstaben . 
Vadå , gruppnavigatör ? 
Jag sitter löst till . Carter också . 
De ersätter oss så snart de hittar några som kan ersätta oss . 
Det lär de inte göra . 
- Varsågod , Croz . 
- Tack , Knifehead . 
- Hör ni ! För 100:e ! 
- Jag har inte hört det förut . 
Aldrig . - Inte ? Croz , Harding vill träffa dig . 
Titta , Egan . Vad gör han tillbaka så tidigt ? 
De har väl fattat sitt beslut . 
- Påfyllning , Mike ? - Gärna det . 
Ni kan sluta undra , mina herrar . 
Ni förstår alla varför jag kom tillbaka i förtid . 
Jösses . Ett nytt uppdrag . 
Flyger vi varje dag numera ? 
230830 , Brady . 30725 , ge det till Cruikshank . 
- Major ? - Clift ! Har vi 230758 ? 
En viktig sak . Jag förstod inte riktigt vad som ... 
Beklagar , sir , men mekanikerna hinner inte få de två planen ni bad om redo till starttiden . Kan vi få en bild av MPI ? Är bomblastlistan skickad till materielavdelningen ? 
Det är klart . De har allt som behövs . 
- Hallå , Croz . - Vi har en . Vi börjar med en tjänstgörande . Homer . Crosby har just befordrats till gruppnavigatör . 
- Välkommen till aphuset , kapten . 
- Tackar . Spence har era fältorder för navigation . 
Kapten , ta det här till S-2 . Tala om vad ni behöver . 
Men för fan . 
Förlåt . Förlåt . 
Hämta en trasa , va ? 
Jösses . Ingen fara . 
TJÄNSTGÖRANDE Häng med , Croz . - Ingen skada skedd . - Tack . 
Det här är ditt kontor . 
Du har en egen jeep . En extraförmån . Om du behöver nåt mer , så säg till Tripp . Okej ? 
Lycka till , Croz . 
Major ? 
Säkert att jag är rätt man för jobbet ? Nej . 
Ert primära mål är Münster . 
Huvudmålet att slå ut är bangårdarna till järnvägsnätet . 
Målet är beläget strax öster om stadskärnan . 
Tystnad . Lyssna nu . 
Så träffsäkerhet är avgörande på det här uppdraget . 
Enligt underrättelser huserar de flesta närbelägna bostäderna järnvägsarbetare . Så om de blir träffade , slår vi ut manskapet som håller de tyska järnvägarna igång . 
Lyse . Överste ? 
Tack , Red . 
95:e i täten med oss lågt , och 390:e överst . 
Det positiva är att det är en kort resa . Münster ligger jäkligt nära . Det positiva är att det är en kort resa . Münster ligger jäkligt nära . 
Det negativa är att vi bara kan få ihop 17 bombplan , varav några inte ens var våra för två dagar sen . Bara 17 bombplan ? 
Det är uppdraget , pojkar : Förstöra transportmöjligheterna för industrin i Ruhr-dalen . Förstått ? 
Ja , sir . 
Bra . Major Egan är befälspilot i Bradys plan . 
Vi har flugit två uppdrag på två dagar . 
Ska man inte rotera skvadronerna ? Så att några får vila ? 
Vilka andra har de ? 
Det är fel . Det är söndag . 
Ja , och imorgon är det måndag . 
Du såg hur nära målpunkten katedralen ligger . 
Vi bombar precis när alla kommer ut ur kyrkan . 
Och ? Det är mycket folk i katedralen . Och i hemmen . 
Och inte bara järnvägsarbetare . 
Alla är delaktiga . 
Vi har aldrig bombat så nära en stads ... Men för tusan , Crank . Det är krig . 
Vårt jobb är att fälla bomber . 
På kvinnor och barn ? 
Kriget slutar inte förrän tyskarna får lida ordentligt . 
Helst innan varenda jäkla kille vi har delat barack med är död eller saknad i strid . 
Ingen av dem vi ska bomba idag sköt ner Buck . 
Tänker du flyga idag eller inte ? 
" Ja , sir . " 
Ja , sir . 
Du ser eländig ut . 
Jag känner mig dålig . Jag tar den . 
Gå och lägg dig , vetja . 
Jag vill se till att alla navigatörer har vad de behöver . 
Jag skulle föredra tyskarnas ovillkorliga kapitulation , men det här duger . Jag skulle föredra tyskarnas ovillkorliga kapitulation , men det här duger . 
Grattis till befordran . 
Gå inte och tro att jag är sur för det . 
Du är ändå den bästa navigatören . 
Du verkar vara ensam om den åsikten . 
Önska mig lycka till i She ' s Gonna . 
She ' s Gonna vadå ? 
Det skulle du vilja veta . 
Hallå ! Stanna lastbilen ! 
- Allt väl , Bucky ? 
- Jadå , fortsätt ni . Jag tar en jeep . 
Jack ! 
- Vi måste byta jacka . - Va ? 
Kom igen . Får jag din jacka . 
Skojar du ? 
Sa de när vi får tillbaka planet ? Inte än . 
Vad heter planet som vi har tilldelats ? 
Royal Flush . 
" Aw-R-Go " ? Vad tusan betyder det ? " Aw-R-Go " ? Vad tusan betyder det ? 
Vi fick det från Framlingham igår . 
Men det flyger . Åtminstone så långt . 
Nu känner jag mig lugnare . 
Tack , Lloyd . 
Har du bytt flygarjacka , major ? 
Buck har jämt avskytt den jackan . 
Den svåraste delen med varje uppdrag var tiden före . Väntan . 
Oavsett hur väl jag plottade rutterna eller hur noggrant jag informerade de andra navigatörerna var jag maktlös när planen väl hade lyft . 
Flanagan lämnar formationen . 
Fan också , en till . 
Befälspilot till akterskytt , ser du vad som är fel med Flanagans plan ? 
Ja , jag ser . Fjärde motorn verkar hacka . 
Stephen tar hans plats i formationen . 
Befälspilot till navigatören , logga det som ännu ett mekaniskt fel . 
Så , har vi mist tre eller fyra plan ? Jag har tappat räkningen . Kom . Så , har vi mist tre eller fyra plan ? Jag har tappat räkningen . 
Kom . Fyra , major . Så vi har 13 plan kvar . 
Fan också ! 
Vi lär inte hinna täta luckan mellan oss och 95:e före kusten . 
Ja , vi ger full kräm . 
Befälspilot till akterskytt , hur långt efter är 390:e ? 
Minst åtta km , sir . 
Tillräckligt stor lucka för att tyskarna ska kunna anfalla oss enskilt . Ja . 
Du , Johnny , det kanske är dags att gå ner och bemanna den tredje kulsprutan , va ? 
Jag är på väg , major . 
Skönt att bli av med honom . 
Han är min andrepilot . 
Han ser bara till att du inte spränger mitt plan . 
Det lär inte ske idag . 
Kulsprutetorn till bombfällare . Klart bombfällaren . 
Är det okej att dra säkringarna ? 
Det är grönt ljus . 
Och syrgas ? Hur är det där bak ? Syrgasen är okej . 
Håll bara patronmatningen redo . Tryck ner matningsreglaget . Håll bara patronmatningen redo . 
Tryck ner matningsreglaget . Matningen är klar . Resten går till skottet . 
Okej , kolla kulsprutorna . - Kulsprutorna klara . - Allt okej ? 
Ja . Kulsprutorna är klara . 
.50-kulsprutorna är klara . 
Jösses . Hur mycket kaffe drack du i morse ? 
Åt helvete för mycket . 
Bomber fällda ! 
Okej , pojkar , jag går ner . Okej . 
Eskortplanen har bränslebrist . De återvänder hem . 
De fick oss över kanalen i alla fall . 
Kulsprutetorn till besättning . Luftvärnseld rakt fram . 
Uppfattat . 
Kulsprutetorn till besättning . Luftvärnseld klockan ett lågt . 
Luftvärnseld klockan tre . Klockan sex . 
Hörru ! - Har jag sagt att jag hatar luftvärnseld ? 
- Inte idag . 
Lauro är träffad . De hoppar . - Fasen . - Jag ser fallskärmar . 
Helvete ! Stymie är nedskjuten . 
Vi är elva kvar . 
Navigatör till befälspilot , tre minuter till referensplatsen . Pilot till navigatör . Uppfattat . 
Harry ? Harry ! 
Nej . - Är vi träffade ? - Harry ! 
Befälspilot till besättning , allt väl där bak ? Kom . 
Clanton ... Halva ansiktet är bortskjutet . 
Jösses . 
För tusan . Harry , andas , Harry . 
Andas . Andas , för tusan ! 
Harry , du får inte dö . 
Andas . 
Snälla , Harry . 
Motor ett lägger av . 
Helvete ! Stäng av bränslet och flöjla den . 
Clanton är död . 
Navigatör till pilot , vi är över referenspunkten . Gira till 057 . 
Uppfattat . Girar till 057 . Kom . 
Luftvärnselden avtar , pojkar . Håll skarp utkik . Det är nog jaktplan överallt . 
Gode Gud . 
Jaktplan klockan tolv . De måste vara hundratals . 
Öppna eld , ge dem vad de tål ! 
Vi förbättrar oddsen . 
Jag är träffad ! 
Jag är träffad i benet ! 
- Mitt ben ! 
- Jag kommer ! 
Pilot till bombfällare , vi närmar oss målet . Är du redo ? Bombfällare till pilot . Svar ja . Pilot till bombfällare . Ta över . Uppfattat . Öppnar bombluckorna . 
Fiendeplan klockan nio högt ! 
Akterskytt . Vi har mist ett till ! Den sista av låga roten . 
Fan också ! 
Motor tre brinner ! 
Stänger av bränslet , och flöjlar . 
Ingen fara ! 
Vi bibehåller hastigheten . Vi bibehåller hastigheten . 
Nätt och jämnt . 
Vi tar oss till målet . 
Cirka en minut till bombfällning . 
Raketer klockan två ! 
Befälspilot till nospartiet . Hur är det där nere ? Vi har bomber att fälla . 
Hambone ! Hambone ! 
De ger sig på oss en gång till . 
Låt det kosta dem dyrt ! 
Jösses , motor fyra stannar ! Vi har bara en motor . 
Hambone är illa sårad . 
Motor två lägger av . Planet skevar redan . Det blir svårt att hålla oss vågrätt . 
- Vi måste lämna formationen . - Helvete . Helvete ! 
Fäll bomberna nu för fan ! 
Larma " överge plan " ! 
Fäll bomberna ! 
Vi ska hoppa ! Fäll bomberna för fan ! 
Förstör bombsiktet ! Skjut sönder det ! 
Jag kan inte hålla planet stadigt länge till ! 
Håll ut , Hambone ! 
Hjälp mig ! Ta hit min fallskärm ! 
Pilot till navigatör , notera i loggen : Skvadronsledaren Egan lämnar formationen . 
Uppfattat . Cruikshank intar ledarposition . 
Uppfattat . Navigatör till pilot , major Egan sjunker snabbt . 
De tänker visst hoppa . 
Kom igen ! Vi måste fort ut ur planet ! 
Hallå , ge mig ett handtag ! 
Petros , sätt fart ! 
Han borde begravas . 
Vi måste få ner Harry . 
George , kom igen , för fan ! Han är död ! George , kom igen , för fan ! Han är död ! Vi måste hoppa ! Kom igen ! 
- Hjälp ! Selen har fastnat ! - Hambone ! 
Hjälp mig loss ! 
Dra i utlösningsmekanismen ! 
De har hoppat ! Allihop ! Nu lämnar vi det här skrället ! 
- Hoppa ! 
- Du först ! - Hoppa ! - Du först ! 
För fan , Brady , jag är din överordnade . Hoppa ! Det är mitt plan ! Du först ! 
Vad fan ! 
Okej . Vi ses , John ! 
Jag är kvar än , era jävlar ! 
Vi är över målet . Släpp bomberna för fan , så vi kan sticka härifrån . 
Bombfällare till pilot . Nu ? Inte före ledarplanet . 
Nu ? 
Vänta . 
Nu ? 
Inte än . 
- Nu . 
- Bomber fällda . 
Där faller de . 
Mitt i prick . 
Inkommande luftvärnseld . 
Hur är det ? 
- Ingen fara med mig . - Vänster midjeskytt till pilot . DeBlasio är träffad i aktern . 
Han blöder , men det är nog ingen fara . 
Uppfattat . 
Pilot till besättning . Luftvärnselden har slutat . Håll utkik . 
Jaktplan klockan tio högt och klockan två högt . 
De ger sig på Cruikshank som ledare . 
Ledarplanet störtar ! 
Jag ser fallskärmar ! 
110:orna är nu klockan fem högt , mot vågrätt . 
Raketer inkommande . Styrbord . 
Jösses , det är hål i vingen ! 
She ' s Gonna är sönderskjutet ! 
Några fallskärmar ? 
Jösses , vi miste just ledarplanet och She ' s Gonna . 
Akterskytt , kulspruteskytt , några fallskärmar ? Jag ser inga . 
Var är alla ? 
Pilot till besättning , ser nån några andra plan från 100:e ? 
- Övre kulspruteskytt , svar nej . 
- Vänster midjeskytt , svar nej . 
Nedre kulspruteskytt , svar nej . 
- Nospartiet , svar nej . - Aktern till pilot , svar nej . - Nospartiet , svar nej . - Aktern till pilot , svar nej . 
Höger midjeskytt , svar nej . 
Fiendeplan klockan fem högt . 
Fler av de jävlarna klockan sju högt . 
Pilot till besättning . Håll i , allihop . 
- Två till kommer . - Klockan två . 
De kommer rakt mot oss . 
Alla kulsprutor redo babord . 
Brassa på , pojkar . 
Håll i , pojkar . Håll i , pojkar . 
Bra skjutet , Milburn . 
Håll skarp utkik , pojkar . De har inte gett upp än . 
Två kommer bakifrån , klockan sex lågt . 
Okej , vänta lite . Jag ska ge dig fritt skottfält . 
Här kommer de , Billy . 
Jag ser dem . Rakt fram . Ta rodret ! 
Klockan tolv vågrätt . 
Vadå ? 
Det är som en klocka . 
Rakt fram är klockan tolv . Så bakom är ... - Klockan sex ? - Just det . 
Öppna eld ! 
Fäll bomberna ! Nu . 
Jag hör dem . 
Inte våra killar . 
Det är 390:e . 
Anropa en av dem via radio . 
Annalkande plan , Station 139 . Bekräfta . 
Plan från 390:e som gör inflygning , detta är tornet . Hör ni mig ? 
Ni har landat på Station 139 . 
Det här är befälhavaren för 100:e . 
Vet ni var min bombgrupp landar ? 
Piloten ? 
Var är våra pojkar , Chick ? 
Ingen av dem klarade sig , sa han . 
Ingen av dem ? 
Här kommer ett till . 
- Det är ett av våra . 
- Vem är det ? 
En av de nya killarna . Rosenthal . 
Det här är plan 087 . Vi har skadade ombord . 
Uppfattat , plan 087 . Vi skickar ut ambulans . 
Var är resten ? 
Gå hem , pojkar . 
- De andra , då ? - Gå hem . 
Kör . 
Lugnt och fint . 
Jag lyfter benen först . 
Vi tar huvudet . 
Försiktigt . 
- Försiktigt . - Vi har honom . 
Vi ska få dig hem , Loren . 
Vad hände med Bubbles ? 
Och Egan ? 
Efter utfrågningen . 
Och Crank ? 
Senare , Kenny . Allihop ? 
Det är nog . 
Det är banne mig nog ! 
Det är sista gången jag går upp . Det är sista gången jag går upp . 
De kan inte tvinga mig . Jag vägrar . 
Jag vägrar . 
Det är banne mig sista gången jag går upp . 
Akternummer 230823 . Invadin ' Maiden . Walts plan . 
Ingen information . Någon ? 
Akternummer 230047 . Sweater Girl . UTFRÅGARE NR 1 Det hör till Atchinsons gäng . 
Ingen information . 
Någon ? 
Akternummer 23534 . Ol ' Dad . 
Ingen information . 
Det var väldigt tufft där uppe , sir . 
Vi hade inte mycket tid för loggar . 
Akternummer 230023 . Forever Yours . Storks besättning . Akternummer 230023 . Forever Yours . Storks besättning . 
Ja , sir . De ... De träffades av en granat . Tidigt . 
Planet brann en stund och sen ... Såg nån några fallskärmar ? 
Akternummer 23229 . Pasadena Nina . 
Ronald ? 
Någon ? 
Akternummer 234423 . She ' s Gonna . 
Bubbles Payne . Navigatör . 
Ingen information . 
Jag såg dem . 
Jaha , vad hände ? 
De brann och sen exploderade de . 
Några fallskärmar ? 
De exploderade , sa jag ju . 
Nej , sir . Inga fallskärmar . 
Akternummer 230087 . Shack Rat . 
Ingen information . 
Akternummer 23237 . Slightly Dangerous . 
Thompsons besättning . 
Ingen information . 
Akternummer 23433 . Leona . 
Ingen information . 
Kära Jean , Du vet redan att din man var den bästa vän jag haft . 
Han var också den bästa navigatör jag nånsin träffat , fast han var för ödmjuk för att medge det för sig själv . fast han var för ödmjuk för att medge det för sig själv . 
Det krävs ett särskilt slags mod för att kunna förbli ödmjuk omgiven av skrytmånsar överallt , men sån var Croz . 
Jag önskar mer än nåt annat att han satt här och inte jag för då behövde ingen skriva det här brevet . 
I NÄSTA AVSNITT Det var ett uppdrag till Münster . Det var ett uppdrag till Münster . Det var tufft . 
Tre uppdrag dina första tre dagar . 
Hundratjugo man dödade på en eftermiddag . 
Jag var inte en av dem . 
Den här miljön är nog inte bra för mig . 
Jag vill återvända till basen . Det här kriget ... Människor ska inte bete sig på det viset . 
När man ser folk förföljas , underkuvas måste man göra nånting . 
Bubbles störtade i förra veckan . Det var mitt fel . 
Gå inte och gråt över det . 
Sätt dig i planet och gör färdigt det jäkla jobbet . 
